hello obj
micro2: Note: Dump of CROM Statements.
width = 72
    constant CROM : CROM_t := (
        --000000000011_111111112222_222222333333_333344444444_445555555555_666666666677_
        --012345678901_234567890123_456789012345_678901234567_890123456789_012345678901_
        b"010010001000_000000000000_000000100001_101101000001_110000000000_111000100000",	-- 0000
        b"100100110000_010000000000_010010100001_101101000001_111001001101_111000100000",	-- 0001
        b"110010000000_000000000000_000110100001_101101000001_000010000001_111000100000",	-- 0002
        b"010010000000_010000000000_000000100001_100001000001_101000010000_111011100000",	-- 0003
        b"010000001000_000111111000_000000100001_111101000001_000000000000_111000000000",	-- 0004
        b"010010001000_000000000000_000000100001_101101000001_000000000001_111000100000",	-- 0005
        b"010010000000_010101111000_000000100001_101101000001_000000000000_111011100000",	-- 0006
        b"010010001000_000110000000_000000100001_101110000000_000000000001_111000100000",	-- 0007
        b"010000001000_000000000000_000000100001_101110000000_111111111110_111000100000",	-- 0010
        b"110001101000_010000000000_000001111101_110011000011_001011000110_111000000000",	-- 0011
        b"010001101000_010000000010_000001101001_110011000010_001011000110_111000000000",	-- 0012
        b"010001101000_010000000010_000001101001_110011000011_001011000110_111000000000",	-- 0013
        b"000110001000_000000000000_001010100001_101110000000_000000000000_111000100000",	-- 0014
        b"011001101000_010000000000_000000100001_101100000000_000000100011_111000000000",	-- 0015
        b"010000001000_000000100000_000000100001_101110000000_111111011011_111000100000",	-- 0016
        b"010111001111_111000000000_000011101001_110011000010_001011000110_111000000000",	-- 0017
        b"100101101000_010000000001_010011101001_110011000010_001011000110_111000000000",	-- 0020
        b"010001101000_110000100010_000001101001_110011000010_001011000110_111000000000",	-- 0021
        b"110010000000_000000000000_000000100001_101001000000_000000001111_111000000000",	-- 0022
        b"010111001111_111000000000_000011101001_110011000011_001011000110_111000000000",	-- 0023
        b"100101101000_010000000001_010011111101_110011000011_001011000110_111000000000",	-- 0024
        b"110000110111_111000000000_000001101001_110011000011_001011000110_111000000000",	-- 0025
        b"010001101000_110000100010_000001101001_110011000011_001011000110_111000000000",	-- 0026
        b"010010001000_000110000000_000000100001_101110000000_000000000010_111000100000",	-- 0027
        b"010010001000_000000100000_000000100001_101110000000_000011111111_111000100000",	-- 0030
        b"000101101000_110000000001_010010100001_111100000000_000000000010_111000000000",	-- 0031
        b"000101101000_010000000001_010010000001_011001000000_000000011010_111000000000",	-- 0032
        b"000101101000_010000000001_010010000100_111100000000_000000000010_111000000000",	-- 0033
        b"000101101000_010000000001_010010000001_011001000000_000000011100_111000000000",	-- 0034
        b"110010000000_000000000000_000000000100_001110000000_000000000000_111000000000",	-- 0035
        b"010010000000_000000000000_000000000011_101100000000_000000000011_111011000000",	-- 0036
        b"100101101000_010000000001_010010100001_111001000000_000000011111_111000000000",	-- 0037
        b"010010001000_000001000000_000000100001_101110000000_000000001111_111000100000",	-- 0040
        b"011111000001_010000000000_000001000001_101100000000_000000000011_111011000000",	-- 0041
        b"101101101000_010000000001_010010100001_111001000000_000000100010_111000000000",	-- 0042
        b"010011000001_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0043
        b"010011111000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0044
        b"110010110000_010000100000_000001101001_110011000011_001011000110_111000000000",	-- 0045
        b"010010001000_000000000000_000000101101_110001000010_001010110011_111000000000",	-- 0046
        b"010000110000_010000000000_000000110101_110001000010_001010110011_111000000000",	-- 0047
        b"010000110000_010000000000_000000111101_110001000010_001010110011_111000000000",	-- 0050
        b"010000110000_010000000000_000000101001_110001000010_001010110011_111000000000",	-- 0051
        b"010000110000_010000000000_000001001101_110001000010_001010110011_111000000000",	-- 0052
        b"010000110000_010000000000_000001010101_110001000010_001010110011_111000000000",	-- 0053
        b"010000110000_010000000000_000001011101_110001000010_001010110011_111000000000",	-- 0054
        b"010000110000_010000000000_000001001001_110001000010_001010110011_111000000000",	-- 0055
        b"110010110000_010000100000_000001101001_110011000011_001011000110_111000000000",	-- 0056
        b"010000110111_111000100000_000001111101_110011000011_000000011001_111000000000",	-- 0057
        b"010010001000_000110000000_000000100001_101110000000_000000000011_111000100000",	-- 0060
        b"010010001000_000000100000_000000100001_101110000000_000001111111_111000100000",	-- 0061
        b"011101101000_110001000000_000000100001_101110000000_000001000000_111000100000",	-- 0062
        b"110111001001_010000000000_010001101001_110001000011_001010110010_111000000000",	-- 0063
        b"110111001001_010000000000_100001101001_110001000011_010011010010_111000000000",	-- 0064
        b"110111001001_010000000000_110001101001_110001000011_011011001101_111000000000",	-- 0065
        b"110111001001_010000000001_000001101001_110001000011_001010110001_111000000000",	-- 0066
        b"110111001001_010000000001_010001101001_110001000011_001010101110_111000000000",	-- 0067
        b"110111001001_010000000001_100001101001_110001000011_001010110000_111000000000",	-- 0070
        b"110111001001_010000000001_110001101001_110001000011_001010101111_111000000000",	-- 0071
        b"010010001000_000000000000_000000100001_110001011100_001010110011_111000000000",	-- 0072
        b"100101101000_010000000000_010010100001_110001011110_001010110011_111000000000",	-- 0073
        b"100101101000_010000000000_010010100001_110001100000_001010110011_111000000000",	-- 0074
        b"100101101000_010000000000_010010100001_110001100010_001010110011_111000000000",	-- 0075
        b"100101101000_010000000000_010010100001_110001100100_001010110011_111000000000",	-- 0076
        b"100101101000_010000000000_010010100001_110001100110_001010110011_111000000000",	-- 0077
        b"100101101000_010000000000_010010100001_110001110110_001010110011_111000000000",	-- 0100
        b"110010000000_000000000000_000000100001_100001000001_001010110111_111000000000",	-- 0101
        b"010000110111_111000100000_000001111101_110011000011_000000110010_111000000000",	-- 0102
        b"010010001000_000110000000_000000100001_101110000000_000000000100_111000100000",	-- 0103
        b"010010001000_000000100001_001100100001_101110000000_000000000111_111000100000",	-- 0104
        b"010010001000_000001000000_000000100001_101110000000_000000000111_111000100000",	-- 0105
        b"010010000000_000000000000_110100100001_101110000000_000000000000_111000000000",	-- 0106
        b"010011000001_010000000000_000000100001_110001000001_001010110111_111000000000",	-- 0107
        b"010000110111_111000100001_001101111101_110011000011_000001000110_111000000000",	-- 0110
        b"010010001000_000110000000_000000100001_101110000000_000000000101_111000100000",	-- 0111
        b"010010001000_000000100001_110100100001_101110000000_000011111111_111000100000",	-- 0112
        b"010010001000_000001000000_000000100001_101110000000_000011111111_111000100000",	-- 0113
        b"010010000000_000000000000_111100100001_101110000000_000000000000_111000000000",	-- 0114
        b"010011000001_010000000000_000000100001_110001000001_001010110111_111000000000",	-- 0115
        b"010000110111_111000100001_110101111101_110011000011_000001001100_111000000000",	-- 0116
        b"110010000000_000000000000_111101111101_100011000011_000001000110_111000000000",	-- 0117
        b"010010001000_000110000000_000000100001_101110000000_000000000110_111000100000",	-- 0120
        b"010010001000_000000100000_000000100001_101110000000_000011111111_111000100000",	-- 0121
        b"010010001000_000010100000_000100100001_101110000000_111111111111_111000100000",	-- 0122
        b"110001101000_110000000001_110100100001_111110000000_000000000000_111000000000",	-- 0123
        b"010010001000_000000000000_000000100001_101110000000_000011111111_111000100000",	-- 0124
        b"000101101000_010001000000_000010100001_111110000000_000000000000_111100000000",	-- 0125
        b"010010001000_000001100000_000000100001_101110000000_000000000111_111000100000",	-- 0126
        b"011001101001_110000000000_000000100001_100011010000_000001100001_111000000000",	-- 0127
        b"110001101001_110000000010_000000100001_111110000000_000000000000_111000100000",	-- 0130
        b"110010000000_000000000000_101100100001_100011111101_000001011100_111000000000",	-- 0131
        b"010010000000_000001100000_110100100001_101110000000_000000000000_111000000000",	-- 0132
        b"110011001001_110000000000_000000100001_111110000000_000000000000_111000100000",	-- 0133
        b"000110001000_000001100000_001010100001_110011000001_000001011110_111000000000",	-- 0134
        b"100101101001_110001100001_010010100001_111110000000_000000000000_111000000000",	-- 0135
        b"110010001000_000000000001_001100100001_111001000000_000001011101_111000000000",	-- 0136
        b"010010010001_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 0137
        b"010010010001_110001000000_000000100001_111110000000_000000000000_111100000000",	-- 0140
        b"010000110111_111010100000_000000100001_111110000000_000000000000_111000000000",	-- 0141
        b"110010000000_000000000000_000001111101_100011000011_000001010110_111000000000",	-- 0142
        b"110010000000_000000000000_000000100001_100001000001_001010110111_111000000000",	-- 0143
        b"010000110111_111000100000_000001111101_110011000011_000001010010_111000000000",	-- 0144
        b"110010000000_000000000000_000110100001_101110000000_000010000001_111000100000",	-- 0145
        b"010010000000_000011100000_000000100001_101110000000_000000000000_111010000000",	-- 0146
        b"010010001000_000110000000_000000100001_101110000000_000000000111_111000100000",	-- 0147
        b"110010000000_000000000000_000000100001_100001000001_001010110100_111000000000",	-- 0150
        b"010010001000_000000100000_000000100001_101110000000_000000000001_111000100000",	-- 0151
        b"110011000111_111000100000_000000100001_010001000001_001010110110_111010000000",	-- 0152
        b"100101101000_110000100000_010011001001_110011000011_000001101010_111000000000",	-- 0153
        b"110011001111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 0154
        b"011000111111_111000000000_000111111101_110011000011_000001101001_111000000000",	-- 0155
        b"010010001000_000110000000_000000100001_101110000000_000000001000_111000100000",	-- 0156
        b"110010000000_000000000000_000000100001_100001000001_001010110100_111000000000",	-- 0157
        b"010011001111_111000100000_000110100001_110001000001_001010110110_111000000000",	-- 0160
        b"011000111111_111000000000_000111111101_110011000011_000001110000_111000000000",	-- 0161
        b"010010001000_000110000000_000000100001_101110000000_000000001001_111000100000",	-- 0162
        b"010010001000_000000100000_101000100001_101110000000_001100111111_111000100000",	-- 0163
        b"010010001000_000001000000_000000100001_101110000000_000000000000_111000100000",	-- 0164
        b"110000001000_000000000001_111110100001_110001000001_001010100111_111000000000",	-- 0165
        b"010010001000_000000100000_100000100001_101110000000_001000000000_111000100000",	-- 0166
        b"010010001000_000001000000_000000100001_101110000000_000000001110_111000100000",	-- 0167
        b"110010001000_000000000001_111110100001_110001000001_001010100111_111100000000",	-- 0170
        b"010010001000_000000000000_000000100001_101110000000_000111000001_111000100000",	-- 0171
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 0172
        b"010010001000_000000000000_000000100001_101110000000_000110000001_111000100000",	-- 0173
        b"110001101000_010000000000_110110100001_110001000001_001010110110_111100100000",	-- 0174
        b"010010001000_000000100000_000000100001_101110000000_000110000000_111000100000",	-- 0175
        b"110010001000_000000000000_100110100001_110001000001_001010110110_111000000000",	-- 0176
        b"110010000000_000000000000_101110100001_101110000000_000000100000_111000000000",	-- 0177
        b"110010000000_000000000000_000000100001_100001000001_001010110110_111000000000",	-- 0200
        b"010010001000_000000100000_000000100001_101110000000_000110001110_111000100000",	-- 0201
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 0202
        b"110010000000_000000000000_000000100001_100001000001_001010110110_111000000000",	-- 0203
        b"110010000000_000000000000_000000100001_100001000001_001010110100_111000000000",	-- 0204
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0205
        b"011000111111_111000000000_000111111101_110011000011_000010000101_111000000000",	-- 0206
        b"010010001000_000010100000_000000100001_101110000000_000010000000_111000100000",	-- 0207
        b"010010001000_000110000000_000000100001_101110000000_000000001010_111000100000",	-- 0210
        b"010001101010_110110001000_000000100001_111110000000_000000000000_111000000000",	-- 0211
        b"010010001000_000001100000_000000100001_101110000000_000011101111_111000100000",	-- 0212
        b"010010001000_000001000000_000000100001_101110000000_000011111111_111000100000",	-- 0213
        b"010010001000_000000000000_000000100001_101110000000_000000011000_111000100000",	-- 0214
        b"010001101001_010000100000_000000100001_110001000001_011111001101_111000000000",	-- 0215
        b"110010000000_000000000000_000000100001_100001000001_011111001001_111000000000",	-- 0216
        b"010011000001_110000100000_000000100001_111110000000_000000000000_111000000000",	-- 0217
        b"010011000001_110000000000_000000100001_110001000001_001010110111_111000000000",	-- 0220
        b"010000110111_111001000000_000001111101_110011000011_000010001100_111000000000",	-- 0221
        b"010010001000_000110010000_000000100001_101110000000_000000010001_111000100000",	-- 0222
        b"110001101010_110000000010_000110100001_111110000000_000000000000_111000000000",	-- 0223
        b"010010001000_000000000000_000000100001_101110000000_110000000000_111000100000",	-- 0224
        b"100100110000_010000000000_010010100001_101110000000_111111111111_111000100000",	-- 0225
        b"010010000000_010000100000_000000100001_101110000000_000000000000_111011100000",	-- 0226
        b"110011000111_111000100000_000000100001_110001000001_011101000000_111010000000",	-- 0227
        b"010010001000_000000000000_000000100001_101110000000_000000010000_111000100000",	-- 0230
        b"110010000000_000000000000_000000100001_100001000001_011111001010_111000000000",	-- 0231
        b"010010001000_000001000000_000000100001_101110000000_000011111111_111000100000",	-- 0232
        b"011011000001_010000000000_000000100001_101110000000_000000000000_111000000000",	-- 0233
        b"010010000000_000000000000_000000100001_101100000000_000000000011_111001100000",	-- 0234
        b"010010001000_000000100000_000000100001_101110000000_000000111111_111000100000",	-- 0235
        b"010011000000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 0236
        b"100100110000_010000000000_010010100001_111001000000_000010011111_111000000000",	-- 0237
        b"010000111000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0240
        b"110001101010_110000000010_000110100001_110001000001_100000010110_111000000000",	-- 0241
        b"010010000000_000000100000_000000100001_100001000001_001010110111_111010000000",	-- 0242
        b"010000010101_111000100010_000001111101_110011000011_000010010111_111000000000",	-- 0243
        b"010010001000_000000000000_000000100001_101110000000_000000001000_111000100000",	-- 0244
        b"010000110101_111010100000_000000100001_110001000001_100000010110_111000000000",	-- 0245
        b"110011000000_010010100000_000001101001_110011000010_000010001000_111000000000",	-- 0246
        b"110010000000_000000000000_000110100001_101110000000_000010000001_111000100000",	-- 0247
        b"110011000111_111011100000_000000100001_110001000001_000111110100_111010000000",	-- 0250
        b"010010001000_000110000000_000000100001_101110000000_000000001011_111000100000",	-- 0251
        b"011110001000_000000000000_000000100001_111110000000_000000000000_111000000000",	-- 0252
        b"010010001000_000000100000_000000100001_101110000000_000111111111_111000100000",	-- 0253
        b"010010000000_110001000000_000000100001_101100000000_000000000011_111011100000",	-- 0254
        b"100100110001_010001000000_010010100001_111001000000_000010101101_111000000000",	-- 0255
        b"100101101001_010001000000_010010100001_111110000000_000000000000_111100100000",	-- 0256
        b"011100111000_010000000000_000000100001_100110000000_100000000000_111000100000",	-- 0257
        b"011100111000_010000000000_000000100001_100110000000_100100000000_111000100000",	-- 0260
        b"011100111000_010000000000_000000100001_100110000000_101000000000_111000100000",	-- 0261
        b"011100111000_010000000000_000000100001_100110000000_101100000000_111000100000",	-- 0262
        b"011100111000_010000000000_000000100001_100110000000_110000000000_111000100000",	-- 0263
        b"011100111000_010000000000_000000100001_100110000000_110100000000_111000100000",	-- 0264
        b"011100111000_010000000000_000000100001_100110000000_111000000000_111000100000",	-- 0265
        b"011100111000_010000000000_000000100001_100110000000_111100000000_111000100000",	-- 0266
        b"010000110111_111000100000_000001111101_110011000011_000010101100_111000000000",	-- 0267
        b"010000111000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0270
        b"010010001000_000001000000_000000100001_101110000000_111111111111_111000100000",	-- 0271
        b"010010001000_000000100000_000000100001_101110000000_000001000101_111000100000",	-- 0272
        b"010011000001_010000000000_000000100001_110001000001_001010110111_111000000000",	-- 0273
        b"010010001000_000110100000_000000100001_101110000000_000000111111_111000100000",	-- 0274
        b"010010001000_000111000001_000000100001_101110000000_000111111111_111000100000",	-- 0275
        b"010010001000_000011111000_000000100001_101110000000_000000010111_111000100000",	-- 0276
        b"010010001000_000111110000_000000100001_111110000000_000000000000_111000000000",	-- 0277
        b"010010001000_000110011000_000000100001_101110000000_000000000011_111000100000",	-- 0300
        b"010000001000_000111101000_000000100001_110100000001_000000000010_111000000000",	-- 0301
        b"000101101110_011110011001_010010100001_111000000000_000000000000_111000000000",	-- 0302
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 0303
        b"010010000000_010101111000_000000100001_101110000000_000000000000_111011100000",	-- 0304
        b"000101101101_111000000001_010010100001_101110000000_111111111111_111000100000",	-- 0305
        b"010010000000_010111011000_000000100001_101110000000_000000000000_111011100000",	-- 0306
        b"010010001000_000000000000_000000100001_101110000000_000000100000_111000100000",	-- 0307
        b"010010000000_010101011000_000000100001_101110000000_000000000000_111011100000",	-- 0310
        b"010010001000_000000000000_000000100001_101110000000_000000000000_111000100000",	-- 0311
        b"011000110000_010111111000_000000100001_101100000000_000000111111_111000000000",	-- 0312
        b"010010001000_000000000000_000000100001_111110000000_000000000000_111000000000",	-- 0313
        b"110010000000_000000000000_000000100001_100001000001_001010100110_111000000000",	-- 0314
        b"100101101000_010000000000_011010100001_111001000000_000011001100_111000000000",	-- 0315
        b"000110001000_000000000000_001010100001_111110000000_000000000000_111000000000",	-- 0316
        b"110010000000_000000000000_000000100001_100001000001_001010100110_111000000000",	-- 0317
        b"000101101000_010000000000_000011101001_110011000011_000011001111_111000000000",	-- 0320
        b"110010000000_000000000000_000110100001_101110000000_000001100101_111000100000",	-- 0321
        b"010010001000_000000000000_000000100001_101110000000_100011100000_111000100000",	-- 0322
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 0323
        b"100100110000_010000000000_010010100001_111100000000_000000000101_111010000000",	-- 0324
        b"110010000000_000000000000_000110100001_101110000000_000001010100_111000100000",	-- 0325
        b"010010001000_000010000000_000000100001_101110000000_000000000111_111000100000",	-- 0326
        b"010010000000_000001100000_000000100001_101100000000_000000000001_111010000000",	-- 0327
        b"010010001000_000000000000_000000100001_101110000000_110101100000_111000100000",	-- 0330
        b"100100110000_010000000000_010010100001_111001000000_000011011001_111000000000",	-- 0331
        b"011000110001_110010000000_001010100001_111110000000_000000000000_100001000000",	-- 0332
        b"010001101000_010000000000_001010100001_011110000000_000000000000_101001000000",	-- 0333
        b"010000110111_111010000000_000001111101_110011000011_000011011010_111000000000",	-- 0334
        b"110010000000_000000000000_000110100001_101110000000_000001000100_111000100000",	-- 0335
        b"010010000000_000100111000_000000100001_101110000000_000000000000_111010000000",	-- 0336
        b"110010000000_000000000000_000110100001_101110000000_000000011110_111000100000",	-- 0337
        b"010010000000_000110111000_000000100001_100001000001_001001111100_111010000000",	-- 0340
        b"110010000000_000000000000_000000100001_100001000001_000101110111_111000000000",	-- 0341
        b"110010000000_000000000000_000000100001_101011100010_000011100111_111000000000",	-- 0342
        b"110010000000_000000000000_000000100001_100001010001_100001101100_111000000000",	-- 0343
        b"110010000000_000000000000_000110100001_101110000000_000001110011_111000100000",	-- 0344
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 0345
        b"010001101000_010000000000_000001101001_110011000011_000000000000_111000100000",	-- 0346
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0347
        b"010010000000_000000000000_000001101001_100011000010_000011101011_111010000000",	-- 0350
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 0351
        b"010010000000_000000100000_000001101001_100011000010_000011111010_111010000000",	-- 0352
        b"110010000000_000000000000_000000100001_101011100010_001100010000_111000000000",	-- 0353
        b"110010000000_000000000000_000000100001_100001000001_000011101110_111000000000",	-- 0354
        b"110010000000_000000000000_000000100001_101011000001_000011100010_111000000000",	-- 0355
        b"110010000000_000000000000_000110100001_101110000000_000101110011_111000100000",	-- 0356
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 0357
        b"010010000000_000000000000_111100100001_101110000000_000000000000_111000000000",	-- 0360
        b"010010000000_000000000000_110100100001_101110000000_000000000000_111000000000",	-- 0361
        b"010010001000_000010100000_000000100001_101110000000_000010000000_111000100000",	-- 0362
        b"110010000000_000000000000_000000100001_100001000001_011111001001_111000000000",	-- 0363
        b"010001101000_010000000000_000000100001_110001000001_011111000111_111000000000",	-- 0364
        b"010001101000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0365
        b"010010001000_000000000000_000000100001_101110000000_000000010000_111000100000",	-- 0366
        b"110010000000_000000000000_000000100001_100001000001_011111001010_111000000000",	-- 0367
        b"010001101000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 0370
        b"010010000000_000000000000_000000100001_101010000001_000000000000_111001100000",	-- 0371
        b"010010001000_000010000000_000000100001_110001000001_000101001100_111000000000",	-- 0372
        b"010010001000_000000100000_000000100001_101110000000_000000001101_111000100000",	-- 0373
        b"110000100000_010000100000_000001101001_110011000010_000101000101_111000000000",	-- 0374
        b"010010001000_000000100000_000000100001_101110000000_000000101100_111000100000",	-- 0375
        b"110000100000_010000100000_000001101001_110011000010_000101001001_111000000000",	-- 0376
        b"110010000000_000000000000_000000100001_100011000001_000100001001_111000000000",	-- 0377
        b"110010000000_000000000000_000000100001_100001000001_001000000100_111000000000",	-- 0400
        b"010010001000_000000100000_000000100001_101110000000_000000100000_111000100000",	-- 0401
        b"110000100000_110000000000_000001101001_110011000010_000100010000_111000000000",	-- 0402
        b"010010001000_000000100000_000000100001_101110000000_000000001101_111000100000",	-- 0403
        b"110000100000_110000000000_000001101001_110011000010_000100010000_111000000000",	-- 0404
        b"010010001000_000000100000_000000100001_101110000000_000000101100_111000100000",	-- 0405
        b"110000100000_110000000000_000001101001_110011000010_000100010000_111000000000",	-- 0406
        b"100101101010_010010000000_010010100001_111100000000_000000000010_111000000000",	-- 0407
        b"100100110010_010010000000_010010100001_111001000000_000100001000_111000000000",	-- 0410
        b"010010001000_000000100000_000000100001_101110000000_000001100000_111000100000",	-- 0411
        b"110000100000_010000100000_000001111101_110011000010_000100001111_111000000000",	-- 0412
        b"010010001000_000000100000_000000100001_101110000000_000001111011_111000100000",	-- 0413
        b"110000100000_010000100000_000001111101_110011000011_000100001111_111000000000",	-- 0414
        b"010010001000_000000100000_000000100001_101110000000_000000100000_111000100000",	-- 0415
        b"010010110000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 0416
        b"010000110000_010010000000_000000100001_110011000001_000100000000_111000000000",	-- 0417
        b"110010000000_000000000000_000000100001_100001000001_001000010111_111000000000",	-- 0420
        b"010010001000_000000000000_000000100001_101101000001_000100111111_111000100000",	-- 0421
        b"110010000000_000000000000_000000100001_100001000001_101000001110_111000000000",	-- 0422
        b"010010001000_000000000000_000000100001_101101000001_000001000010_111000100000",	-- 0423
        b"011000100000_010010000010_000001101001_110011000010_001000100110_111000000000",	-- 0424
        b"110000111111_111000000000_000001101001_110011000010_001000011111_111000000000",	-- 0425
        b"011001101000_000000000010_000001101001_110011000010_001000101000_111000000000",	-- 0426
        b"011001101000_000000000010_000001101001_110011000010_001000110010_111000000000",	-- 0427
        b"011001101000_000000000010_000001101001_110011000010_001001000111_111000000000",	-- 0430
        b"010010001000_000000000000_000000100001_101110000000_000001001000_111000100000",	-- 0431
        b"011000100000_010010000010_000001101001_110011000010_001001110101_111000000000",	-- 0432
        b"011101101000_000000000010_000001101001_110011000010_001001111001_111000000000",	-- 0433
        b"010000000000_000000000010_000001101001_110011000010_001000110111_111000000000",	-- 0434
        b"010010001000_000000000000_000000100001_101110000000_000001010010_111000100000",	-- 0435
        b"011000100000_010010000010_000001101001_110011000010_001010000110_111000000000",	-- 0436
        b"011001101000_000000000010_000001101001_110011000010_001010001111_111000000000",	-- 0437
        b"011001101000_000000000010_000001101001_110011000010_001010100100_111000000000",	-- 0440
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 0441
        b"100100110000_010000000000_010010100001_101110000000_100111001000_111000100000",	-- 0442
        b"011000100000_010010000010_000001101001_110011000010_001010010010_111000000000",	-- 0443
        b"011001101000_000000000010_000001101001_110011000010_001010010101_111000000000",	-- 0444
        b"010001101000_010000000000_000000100001_101110000000_001001001001_111000100000",	-- 0445
        b"110000100000_010010000000_000001101001_110011000010_001001011101_111000000000",	-- 0446
        b"010001101000_010000000000_000000100001_101110000000_001001010010_111000100000",	-- 0447
        b"110000100000_010010000000_000001101001_110011000010_001001100110_111000000000",	-- 0450
        b"010001101000_010000000000_000000100001_101110000000_001001010110_111000100000",	-- 0451
        b"110000100000_010010000000_000001101001_110011000010_001001101101_111000000000",	-- 0452
        b"010001101000_010000000000_000000100001_101110000000_001011001001_111000100000",	-- 0453
        b"110000100000_010010000000_000001101001_110011000010_001001100001_111000000000",	-- 0454
        b"010001101000_010000000000_000000100001_101110000000_001011010110_111000100000",	-- 0455
        b"110000100000_010010000000_000001101001_110011000010_001001110001_111000000000",	-- 0456
        b"010001101000_010000000000_000000100001_101110000000_001011010010_111000100000",	-- 0457
        b"110000100000_010010000000_000001101001_110011000010_001001101001_111000000000",	-- 0460
        b"010001101000_010000000000_000000100001_101110000000_100111001101_111000100000",	-- 0461
        b"110000100000_010010000000_000001101001_110011000010_001010100010_111000000000",	-- 0462
        b"010001101000_010000000000_000000100001_101110000000_110101001101_111000100000",	-- 0463
        b"110000100000_010010000000_000001101001_110011000010_001010111001_111000000000",	-- 0464
        b"110010000000_000000000000_000000100001_100001000001_000111110101_111000000000",	-- 0465
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 0466
        b"110010000000_000000000000_000000100001_101011000001_000101000001_111000000000",	-- 0467
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 0470
        b"110010000000_000000000000_000000100001_101011000001_000101000001_111000000000",	-- 0471
        b"010010001000_000000000000_000000100001_101110000000_000000000100_111000100000",	-- 0472
        b"110010000000_000000000000_000000100001_101011000001_000101000001_111000000000",	-- 0473
        b"110010000000_000000000000_000000100001_100001000001_000101011011_111000000000",	-- 0474
        b"110010000000_000000000000_000000100001_100001000001_000101110101_111000000000",	-- 0475
        b"010001101100_110000000000_000000100001_110011000001_000100111111_111000000000",	-- 0476
        b"110010000000_000000000000_000000100001_100001000001_000101011011_111000000000",	-- 0477
        b"010010001000_000000000000_000000100001_101110000000_000000000101_111000100000",	-- 0500
        b"010010001000_000010100000_000000100001_101110000000_000001000011_111000100000",	-- 0501
        b"010001101000_010010000000_000000100001_110001000001_000101101110_111000000000",	-- 0502
        b"010010000010_010000000000_000000100001_100001000001_000101100000_111011100000",	-- 0503
        b"110010000000_000000000000_000000100001_101011000001_000101000110_111000000000",	-- 0504
        b"110010000000_000000000000_000000100001_100001000001_000111110101_111000000000",	-- 0505
        b"110010000000_000000000000_000110100001_101101000001_000011000000_111000100000",	-- 0506
        b"010010000000_000000000000_000000100001_101101000001_000000000000_111010000000",	-- 0507
        b"110011000100_111000000000_000001101001_110001000010_000101110111_111000000000",	-- 0510
        b"010010001000_000000000000_000000100001_110001000001_001010100000_111000000000",	-- 0511
        b"010010001000_000000000000_000000100001_110001000001_101000001110_111000000000",	-- 0512
        b"110010000000_000000000000_000000100001_101011000001_000011100010_111000000000",	-- 0513
        b"110010000000_000000000000_000000100001_100001000001_001000000100_111000000000",	-- 0514
        b"010010001000_000000100000_000000100001_101110000000_000000100000_111000100000",	-- 0515
        b"110000100000_010000100000_000001101001_110011000010_000101001100_111000000000",	-- 0516
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 0517
        b"010010001000_000010000000_000000010010_110001000001_000101001100_111000000000",	-- 0520
        b"010010001000_000000100000_000000100001_101110000000_000000110111_111000100000",	-- 0521
        b"110000100000_110000000000_000001111101_110011000010_000101011001_111000000000",	-- 0522
        b"010010001000_000000100000_000000100001_101110000000_000000110000_111000100000",	-- 0523
        b"010000010000_110000000010_000001111101_110011000010_000101011001_111000000000",	-- 0524
        b"100100110010_010010000000_010010010000_111110000000_000000000000_111000000000",	-- 0525
        b"100101101010_010010000000_010010100001_111110000000_000000000000_111000000000",	-- 0526
        b"010000110000_010010000000_000000100001_110001000001_001000000100_111000000000",	-- 0527
        b"110010000000_000000000000_000000100001_100011000001_000101010001_111000000000",	-- 0530
        b"110010000000_000000000000_000000100001_100001000001_001000010111_111000000000",	-- 0531
        b"010001101010_010000000000_000000100001_111010000001_000000000000_111000000000",	-- 0532
        b"110010000000_000000000000_000000100001_100001000001_000101100000_111000000000",	-- 0533
        b"010010001000_000000000000_000000100001_101110000000_000000101100_111000100000",	-- 0534
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0535
        b"110010000000_000000000000_000110100001_101110000000_000100101100_111000100000",	-- 0536
        b"010010000000_000000000000_000000100001_100011000001_000101100000_111010000000",	-- 0537
        b"010010001000_000010100000_000000100001_101110000000_000000000110_111000100000",	-- 0540
        b"110010000000_000000000000_000110100001_101110000000_000100101100_111000100000",	-- 0541
        b"110010000000_000000000000_000000100001_101100000000_000000000010_111000000000",	-- 0542
        b"100101101000_010000000001_010010100001_111001000000_000101100011_111010000000",	-- 0543
        b"010010001000_000000100000_000000100001_101110000000_000000000111_111000100000",	-- 0544
        b"011111000000_110000000000_000000100001_101110000000_000000110000_111000100000",	-- 0545
        b"010000111000_010000000000_000000100001_110001000001_000110000111_111000000000",	-- 0546
        b"110010000000_000000000000_000110100001_101110000000_000100101100_111000100000",	-- 0547
        b"010000110111_111010100000_000000100001_011110000000_000000000000_111000000000",	-- 0550
        b"010010000000_000000000000_000001001001_100011000011_000101100010_111010000000",	-- 0551
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 0552
        b"010010001000_000000000000_000000100001_101110000000_000001011110_111000100000",	-- 0553
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0554
        b"010001101010_110000000000_000000100001_110011000001_000110000111_111000000000",	-- 0555
        b"110010000000_000000000000_000000100001_100001000001_000110000100_111000000000",	-- 0556
        b"010010001000_000000000000_000000100001_101110000000_000000011100_111000100000",	-- 0557
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0560
        b"010010001000_000000000000_000000100001_101110000000_000000111111_111000100000",	-- 0561
        b"110010000000_000000000000_000000100001_100011000001_000101101100_111000000000",	-- 0562
        b"010010001000_000000000000_000000100001_101110000000_000000101111_111000100000",	-- 0563
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0564
        b"010010001000_000000000000_000000100001_101110000000_000000100000_111000100000",	-- 0565
        b"110010000000_000000000000_000000100001_100011000001_000110000111_111000000000",	-- 0566
        b"110010000000_000000000000_000000100001_100001000001_000110000100_111000000000",	-- 0567
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0570
        b"010010000000_000000000000_000001101001_101010000011_000000000000_111010000000",	-- 0571
        b"010010001000_000000000000_000000100001_101110000000_000001001011_111000100000",	-- 0572
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0573
        b"010010001000_000000000000_000000100001_101110000000_000001010100_111000100000",	-- 0574
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0575
        b"010010001000_000000000000_000000100001_101110000000_000000110010_111000100000",	-- 0576
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0577
        b"010010001000_000000000000_000000100001_101110000000_000000110000_111000100000",	-- 0600
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0601
        b"010010001000_000000000000_000000100001_101110000000_000000111110_111000100000",	-- 0602
        b"110010000000_000000000000_000000100001_100011000001_000110000111_111000000000",	-- 0603
        b"010010001000_000000000000_000000100001_101110000000_000000001101_111000100000",	-- 0604
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0605
        b"010010001000_000000000000_000000100001_101110000000_000000001010_111000100000",	-- 0606
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 0607
        b"010010001000_000000100000_000000100001_101110000000_000000000001_111000100000",	-- 0610
        b"011101101000_110000100000_000000100001_101110000000_000000000000_111010000000",	-- 0611
        b"110011001000_110000000000_000001101001_111010000011_000000000000_111000000000",	-- 0612
        b"110010000000_000000000000_000110100001_101110000000_000011000010_111000100000",	-- 0613
        b"010010001000_000000100000_000000100001_101110000000_000011011111_111000100000",	-- 0614
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 0615
        b"110000100000_110001000000_000001101001_111010000010_000000000000_111000000000",	-- 0616
        b"110010000000_000000000000_000000100001_100001000001_001000000101_111000000000",	-- 0617
        b"110011000111_111000100000_000000100001_111110000000_000000000000_111010000000",	-- 0620
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 0621
        b"010010000000_000000000000_000001101001_100001000010_000111111111_111010000000",	-- 0622
        b"010010001000_000010101000_000000100001_110011000001_011110111101_111000000000",	-- 0623
        b"010011001111_111000000000_000001101001_111011000010_011110001011_111000000000",	-- 0624
        b"010010001000_000000100000_000000100001_101110000000_000000000011_111000100000",	-- 0625
        b"110000011000_110000000010_000001101001_110011000010_000111010010_111000000000",	-- 0626
        b"010010001000_000000100000_000000100001_101110000000_000000001111_111000100000",	-- 0627
        b"010000010000_010000100010_000001101001_110011000010_000111011100_111000000000",	-- 0630
        b"010000000000_000000100010_000001101001_110011000010_000111110000_111000000000",	-- 0631
        b"010000000000_000000100010_000001101001_110011000010_000111100110_111000000000",	-- 0632
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0633
        b"010010000000_000001000000_000001101001_100011000011_000110110111_111010000000",	-- 0634
        b"110000110000_110111111000_000001101001_110011000010_000111000011_111000000000",	-- 0635
        b"010000000000_000000100010_000001101001_110011000010_000111010010_111000000000",	-- 0636
        b"010010001000_000000100000_000000100001_101110000000_000000011010_111000100000",	-- 0637
        b"110000011000_110000000010_000001101001_110011000010_000111101100_111000000000",	-- 0640
        b"010010001000_000000100000_000000100001_101110000000_000001111111_111000100000",	-- 0641
        b"110000011000_110000000010_000001101001_110011000010_000110111100_111000000000",	-- 0642
        b"110010000000_000000000000_000110100001_101110000000_000011100000_111000100000",	-- 0643
        b"010010001000_000000100000_000000100001_101110000000_000100000111_111000100000",	-- 0644
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 0645
        b"110000100000_110001000000_000001101001_110011000010_000110111001_111000000000",	-- 0646
        b"010010001000_000000100000_000000100001_101110000000_000000001101_111000100000",	-- 0647
        b"110000100000_010000100000_000001101001_110011000010_000110101011_111000000000",	-- 0650
        b"010010001000_000010100000_000000100001_101110000000_000000001010_111000100000",	-- 0651
        b"110000100010_110000000000_000001101001_110011000011_000110110101_111000000000",	-- 0652
        b"010001101000_110000000000_000000100001_110001000001_001000000001_111000000000",	-- 0653
        b"110010000000_000000000000_000000100001_100001000001_000110110011_111000000000",	-- 0654
        b"110010000000_000000000000_000000100001_100001000001_000110000100_111000000000",	-- 0655
        b"110010000000_000000000000_000000100001_101011100011_011110001011_111000000000",	-- 0656
        b"110010000000_000000000000_000110100001_101110000000_000101010000_111000100000",	-- 0657
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0660
        b"010010001000_000000000000_000000100001_110001000001_101000001111_111000000000",	-- 0661
        b"010001101110_010100011001_001100100001_110011000001_000011100111_111000000000",	-- 0662
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0663
        b"110010000000_000000000000_000000100001_100011000001_000111111010_111000000000",	-- 0664
        b"010001101000_010010100000_000000100001_110001000001_001000000001_111000000000",	-- 0665
        b"010001101010_110000000000_000000100001_111011000001_000110111010_111000000000",	-- 0666
        b"110010000000_000000000000_000110100001_101110000000_000011000001_111000100000",	-- 0667
        b"110000001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0670
        b"010010001000_000000000000_000000100001_101110000000_000000000111_111000100000",	-- 0671
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0672
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 0673
        b"011001101111_010000000000_000110100001_101110000000_000011100000_111000100000",	-- 0674
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 0675
        b"011111001000_010000100000_000000100001_101110000000_000011100001_111000100000",	-- 0676
        b"110000100000_110000000000_000001101001_111011000010_011110001011_111000000000",	-- 0677
        b"110010000000_000000000000_000000100001_100001000001_001000011000_111000000000",	-- 0700
        b"010010001000_000000000000_000000100001_101110000000_000001011100_111000100000",	-- 0701
        b"110010000000_000000000000_000000100001_101011000001_000110111010_111000000000",	-- 0702
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 0703
        b"010010000000_000000100000_000001101001_101011000011_011110001011_111010000000",	-- 0704
        b"010010001000_000010100000_000000100001_101110000000_000001010010_111000100000",	-- 0705
        b"110010000000_000000000000_000000100001_100001000001_000101101011_111000000000",	-- 0706
        b"110010000000_000000000000_000000100001_100001000001_000101110111_111000000000",	-- 0707
        b"110010000000_000000000000_000000100001_100001000001_000110110011_111000000000",	-- 0710
        b"110010000000_000000000000_000000100001_100011000001_000111001100_111000000000",	-- 0711
        b"110010000000_000000000000_000000100001_100001000001_001000000100_111000000000",	-- 0712
        b"110010000000_000000000000_000000100001_100001000001_000110000111_111000000000",	-- 0713
        b"110010000000_000000000000_000110100001_101110000000_000011100000_111000100000",	-- 0714
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 0715
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0716
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 0717
        b"110010110000_010000100000_000001101001_110011000011_000111001010_111000000000",	-- 0720
        b"110010001000_000000000000_000000100001_111011000001_011110001011_111010000000",	-- 0721
        b"010010001000_000010100000_000000100001_101110000000_000001000000_111000100000",	-- 0722
        b"010000111010_110010100000_000000100001_110001000001_000111110100_111000000000",	-- 0723
        b"010001101100_111000000000_000000100001_101110000000_000000000011_111000100000",	-- 0724
        b"110010000000_000000000000_000000100001_100001000001_000111100011_111000000000",	-- 0725
        b"110010000000_000000000000_000000100001_100001000001_000101101011_111000000000",	-- 0726
        b"110010000000_000000000000_000000100001_100001000001_000101110111_111000000000",	-- 0727
        b"010010001000_000000000000_000000100001_110001000001_001010100000_111000000000",	-- 0730
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 0731
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 0732
        b"110010000000_000000000000_000000100001_100011000001_000111100011_111000000000",	-- 0733
        b"110010000000_000000000000_000000100001_100001000001_000111111100_111000000000",	-- 0734
        b"010010001000_000010100000_000000100001_101110000000_000001001111_111000100000",	-- 0735
        b"110010000000_000000000000_000000100001_100001000001_000101101011_111000000000",	-- 0736
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 0737
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 0740
        b"011101101000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 0741
        b"110010111000_010000000000_000000100001_111011000001_011110001011_111010000000",	-- 0742
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 0743
        b"011101110000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 0744
        b"110011001000_010000000000_000000100001_111010000001_000000000000_111010000000",	-- 0745
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 0746
        b"110010000000_000000000000_000000100001_100001000001_000111101001_111000000000",	-- 0747
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 0750
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 0751
        b"011101101000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 0752
        b"110011111000_010000000000_000000100001_111010000001_000000000000_111010000000",	-- 0753
        b"110010000000_000000000000_000000100001_101011100011_011110001011_111000000000",	-- 0754
        b"010010001000_000010100000_000000100001_101110000000_000001011010_111000100000",	-- 0755
        b"110010000000_000000000000_000000100001_100001000001_000101101011_111000000000",	-- 0756
        b"010001101100_111000000000_000000100001_110001000001_000111101001_111000000000",	-- 0757
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 0760
        b"110010000000_000000000000_000000100001_100001000001_000111100011_111000000000",	-- 0761
        b"110010000000_000000000000_000000100001_100001000001_011110111101_111000000000",	-- 0762
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 0763
        b"110010000000_000000000000_000000100001_100001000001_000111111100_111000000000",	-- 0764
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 0765
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0766
        b"110010000000_000000000000_000110100001_101110000000_000011000001_111000100000",	-- 0767
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0770
        b"110010000000_000000000000_000110100001_101110000000_000011100000_111000100000",	-- 0771
        b"010010001000_000000000000_000000100001_101110000000_000011100001_111000100000",	-- 0772
        b"110011000111_111000000000_000000100001_111010000001_000000000000_111010000000",	-- 0773
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 0774
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 0775
        b"110010000000_000000000000_000110100001_101110000000_000011000010_111000100000",	-- 0776
        b"010010001000_000000000000_000000100001_101110000000_000011000011_111000100000",	-- 0777
        b"110011000111_111000000000_000000100001_111010000001_000000000000_111010000000",	-- 1000
        b"110010000000_000000000000_000110100001_101110000000_000011100000_111000100000",	-- 1001
        b"110010000000_000000000000_000000100001_100001000001_001000000101_111000000000",	-- 1002
        b"110011000111_111000100000_000000100001_111010000001_000000000000_111010000000",	-- 1003
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 1004
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 1005
        b"010000110111_110000100000_000001111101_110011000011_001000001010_111000000000",	-- 1006
        b"010010001000_000001000000_000000100001_101110000000_000000000100_111000100000",	-- 1007
        b"010010000001_010000101000_000000100001_101110000000_000000000000_111011100000",	-- 1010
        b"010001101000_110000110010_000000100001_111110000000_000000000000_111000000000",	-- 1011
        b"110011000111_111000100000_000110100001_111110000000_000000000000_111010000000",	-- 1012
        b"010010001000_000001000000_000000100001_101110000000_000001001111_111000100000",	-- 1013
        b"011111000001_010000000000_000000100001_100011000001_001000010001_111010000000",	-- 1014
        b"000101101000_010000000000_000010100001_111110000000_000000000000_111000000000",	-- 1015
        b"101101101001_010001000000_110010100001_111100000000_000000000101_111000000000",	-- 1016
        b"000101101000_010000000000_000010100001_111110000000_000000000000_111000000000",	-- 1017
        b"101101101001_010001000000_110010100001_111001000000_001000001111_111000000000",	-- 1020
        b"010000110111_110000100000_000001111101_110011000011_001000001101_111000000000",	-- 1021
        b"010010001000_000000100000_000000100001_101110000000_000001001111_111000100000",	-- 1022
        b"010011000000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 1023
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 1024
        b"010010010001_010000100000_000000100001_111110000000_000000000000_111000000000",	-- 1025
        b"010011111000_110000100000_000000100001_111010000001_000000000000_111000000000",	-- 1026
        b"110010000000_000000000000_000110100001_101110000000_000011100001_111000100000",	-- 1027
        b"010010001000_000000100000_000000100001_101110000000_000000000100_111000100000",	-- 1030
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 1031
        b"011101000000_010000110000_000000100001_101110000000_000000000000_111011100000",	-- 1032
        b"110000101000_110000000010_000000100001_011110000000_000000000000_111000000000",	-- 1033
        b"010000110101_111000000000_000001001001_110011000011_101000010000_111000000000",	-- 1034
        b"010010001000_000000001000_000000100001_111110000000_000000000000_111000000000",	-- 1035
        b"010000110111_111000000000_000000100001_110011000001_101000010000_111000000000",	-- 1036
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1037
        b"110010000000_000000000000_000110100001_101110000000_000100100010_111000100000",	-- 1040
        b"110011000111_111000000000_000000100001_110001000001_000101010000_111010000000",	-- 1041
        b"110010000000_000000000000_000110100001_101110000000_000100100100_111000100000",	-- 1042
        b"110011000111_111000000000_000000100001_110001000001_000101010000_111010000000",	-- 1043
        b"110010000000_000000000000_000110100001_101110000000_000100100011_111000100000",	-- 1044
        b"110011000111_111000000000_000000100001_110011000001_000101001001_111010000000",	-- 1045
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1046
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1047
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1050
        b"110010000000_000000000000_011000100001_100001000001_001000101111_111000000000",	-- 1051
        b"010001101100_111000000000_000000100001_110001000001_000111101001_111000000000",	-- 1052
        b"110010000000_000000000000_000000100001_100001000001_011110111101_111000000000",	-- 1053
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 1054
        b"110010001000_000000000001_001000100001_110001000001_011010001110_111010000000",	-- 1055
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1056
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1057
        b"110010000000_000000000000_000000101001_101010000010_000000000000_111000000000",	-- 1060
        b"010001101000_010011100000_000000100001_111010000001_000000000000_111000000000",	-- 1061
        b"010010001000_000000000000_000000010100_110001000001_001001001101_111000000000",	-- 1062
        b"110010000000_000000000000_000000100001_100001000001_100111000100_111000000000",	-- 1063
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1064
        b"010001101000_010100100000_000000101001_110011000011_001000110011_111000000000",	-- 1065
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1066
        b"110010000000_000000000000_000000100001_100001000001_001000111110_111000000000",	-- 1067
        b"010001101100_110011011000_000000101001_110011000010_001001011000_111000000000",	-- 1070
        b"110010000000_000000000000_000000100001_100001000001_001000111110_111000000000",	-- 1071
        b"110010000000_000000000000_000000101001_100011000010_000101001001_111000000000",	-- 1072
        b"110010000000_000000000000_000110100001_101110000000_000100100101_111000100000",	-- 1073
        b"110001101011_011000000000_000000100001_110001000001_100111000100_111010000000",	-- 1074
        b"010001101011_011011011010_000000100001_110011000001_001000111001_111000000000",	-- 1075
        b"010010001000_000100100000_000000010010_110001000001_000101001100_111000000000",	-- 1076
        b"010010001000_000000100000_000000100001_101110000000_000000111101_111000100000",	-- 1077
        b"110000100000_010000100000_000001111101_110011000010_000101011001_111000000000",	-- 1100
        b"010010001000_000000100000_000000100001_101110000000_000001111101_111000100000",	-- 1101
        b"110000100000_010000100000_000001111101_110011000011_000101011001_111000000000",	-- 1102
        b"010011000110_110000000000_000000100001_111100000000_000000000010_111000000000",	-- 1103
        b"100100110100_110100100000_010010100001_111001000000_001001000100_111000000000",	-- 1104
        b"010000110000_010100100000_000000010000_110001000001_001000000100_111000000000",	-- 1105
        b"110010000000_000000000000_000000100001_100011000001_001000111111_111000000000",	-- 1106
        b"010010001000_000000000000_000000100001_101110000000_001001001001_111000100000",	-- 1107
        b"110010000000_000000000000_000000010110_100001000001_001001001101_111000000000",	-- 1110
        b"010001101011_011011011000_001010100001_111110000000_000000000000_001001000000",	-- 1111
        b"110010000000_000000000000_000000100001_100001000001_100101111011_111000000000",	-- 1112
        b"010001101100_110000000000_000000100001_110001000001_000101011011_111000000000",	-- 1113
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1114
        b"110001101000_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 1115
        b"110010000000_000000000000_000001101001_100001000011_001010100000_111000000000",	-- 1116
        b"010010001000_000000000000_000000100001_101110000000_000100111100_111000100000",	-- 1117
        b"110010000000_000000000000_000000110101_100001000010_101000001110_111000000000",	-- 1120
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1121
        b"110010000000_000000000000_000110100001_101110000000_000100100101_111000100000",	-- 1122
        b"110010000000_000000000000_000000101001_100011000011_001001010101_111000000000",	-- 1123
        b"010010000000_000000000000_000000110101_100011000011_001001011000_111010000000",	-- 1124
        b"010001101000_010100000000_000000110101_110011000010_001001011010_111010000000",	-- 1125
        b"010001101100_010011011000_000000100001_110001000001_000101010000_111000000000",	-- 1126
        b"010001101000_010100100000_000000101001_111010000011_000000000000_111000000000",	-- 1127
        b"010010001000_000000000000_000000100001_101110000000_000000000011_111000100000",	-- 1130
        b"110010000000_000000000000_000000100001_101011000001_000101000001_111000000000",	-- 1131
        b"010001101100_010011011000_000000100001_110001000001_000110000100_111000000000",	-- 1132
        b"010001101011_011000000000_000000100001_110001000001_000101011011_111000000000",	-- 1133
        b"110010000000_000000000000_000000100001_100011000001_000101110011_111000000000",	-- 1134
        b"010010001000_000000000000_000000010100_110001000001_001001001101_111000000000",	-- 1135
        b"010001101000_010101100000_000000100001_110001000001_100000100010_111000000000",	-- 1136
        b"110010000000_000000000000_000000101101_100011000010_000100111010_111000000000",	-- 1137
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1140
        b"010010001000_000000000000_000000010110_110001000001_001001001101_111000000000",	-- 1141
        b"110010000000_000000000000_000000100001_100001000001_001101100000_111000000000",	-- 1142
        b"110010000000_000000000000_000000101101_101011000010_000100111010_111000000000",	-- 1143
        b"010001101101_110000000000_000000100001_110001000001_000101011011_111000000000",	-- 1144
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1145
        b"010010001000_000000000000_000000010100_110001000001_001001001101_111000000000",	-- 1146
        b"110001101011_011000000000_000110100001_111110000000_000000000000_111000000000",	-- 1147
        b"110011000111_111100100000_000000100001_110011000001_000101001001_111010000000",	-- 1150
        b"010010001000_000000000000_000000010110_110001000001_001001001101_111000000000",	-- 1151
        b"110001101011_011000000000_000110100001_111110000000_000000000000_111000000000",	-- 1152
        b"010010000000_000000000000_000000100001_100001000001_000101011011_111010000000",	-- 1153
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1154
        b"010010001000_000000000000_000000100001_101101000001_001001101111_111000100000",	-- 1155
        b"110010000000_000000000000_000000010100_100001000001_001001001101_111000000000",	-- 1156
        b"110010000000_000000000000_010000100001_100001000001_100111001001_111000000000",	-- 1157
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1160
        b"010010001000_000000000000_000000100001_101110000000_001001110011_111000100000",	-- 1161
        b"110010000000_000000000000_000000010110_100001000001_001001001101_111000000000",	-- 1162
        b"110010000000_000000000000_010000100001_100001000001_100110110010_111000000000",	-- 1163
        b"110010000000_000000000000_000000100001_100011000001_001001001011_111000000000",	-- 1164
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 1165
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 1166
        b"110001101110_110000000001_110100100001_111011100011_001011001000_111000000000",	-- 1167
        b"110011000111_111000000001_000000100001_111011000001_001011001000_111010000000",	-- 1170
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1171
        b"110010000000_000000000000_000000100001_100001000001_001001111100_111000000000",	-- 1172
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1173
        b"010010001000_000000011000_100000100001_111110000000_000000000000_111000000000",	-- 1174
        b"010010001000_000001111000_110000100001_111110000000_000000000000_111000000000",	-- 1175
        b"010010001000_000010011000_011000100001_111110000000_000000000000_111000000000",	-- 1176
        b"010010001000_000010111001_100000100001_111110000000_000000000000_111000000000",	-- 1177
        b"110010000000_000000000000_000110100001_101110000000_000000100001_111000100000",	-- 1200
        b"010010000000_000000000001_010000100001_101110000000_000000000000_111010000000",	-- 1201
        b"010001110000_010000000000_000000100001_101110000000_000010000000_111000100000",	-- 1202
        b"110010000000_000000000000_000110100001_101110000000_000101110010_111000100000",	-- 1203
        b"110011000111_111000000001_110000100001_110001000001_011010001000_111010000000",	-- 1204
        b"110010000000_000000000000_000000100001_100011000001_011001001111_111000000000",	-- 1205
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1206
        b"110010000000_000000000000_000110100001_101110000000_000011000001_111000100000",	-- 1207
        b"011001111000_010000000010_000000100001_010001000001_001010001110_111000000000",	-- 1210
        b"110001101000_010000000010_000001101000_110011000010_000101001001_111010000000",	-- 1211
        b"110001101000_010000000000_000001111101_110011000010_001010001100_111000000000",	-- 1212
        b"110011001111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 1213
        b"110010000000_000000000000_000000100001_100001000001_000110110011_111000000000",	-- 1214
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1215
        b"010010000000_000000000000_000000100001_101010000001_000000000000_111010000000",	-- 1216
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1217
        b"110010000000_000000000000_000000100001_100001000001_001001111100_111000000000",	-- 1220
        b"110010000000_000000000000_000000100001_100011000001_001000101000_111000000000",	-- 1221
        b"010010001000_000011011000_000000100001_101110000000_000000011000_111000100000",	-- 1222
        b"010000001000_000100100000_000000100001_110001000001_100111000100_111000000000",	-- 1223
        b"110010000000_000000000000_000000100001_100011000001_000101001001_111000000000",	-- 1224
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1225
        b"110010000000_000000000000_011000100001_100001000001_001000101111_111000000000",	-- 1226
        b"010010001000_000000000000_000000100001_110001000001_101000001110_111000000000",	-- 1227
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 1230
        b"010010001000_000000100000_000000100001_101110000000_000000000011_111000100000",	-- 1231
        b"010010001000_000000000000_000000100001_101110000000_001010011111_111000100000",	-- 1232
        b"110011000111_111000100000_000000100001_110001000001_001010100000_111010000000",	-- 1233
        b"110010000000_000000000000_000000100001_100001000001_011010001110_111000000000",	-- 1234
        b"010010001000_000000000000_000000100001_110001000001_101000001110_111000000000",	-- 1235
        b"011101101011_110100000001_111110100001_111011000001_001100010011_111000000000",	-- 1236
        b"010000110111_111011110000_000000100001_110011000001_001010011110_111000000000",	-- 1237
        b"110010000000_000000000000_000110100001_101110000000_000001110011_111000100000",	-- 1240
        b"110011000111_111000000000_000000100001_111010000001_000000000000_111010000000",	-- 1241
        b"110010000000_000000000000_000000100001_100001000001_000101010000_111000000000",	-- 1242
        b"110001101000_010000000000_000000100001_110011000001_000000000000_111000100000",	-- 1243
        b"110010000000_000000000000_000000100001_100011100010_000100111000_111000000000",	-- 1244
        b"110010000000_000000000000_000000100001_100011000001_000000000100_111000000000",	-- 1245
        b"011001101000_000000000010_000110100001_110011000001_101000010000_111000000000",	-- 1246
        b"110010000000_000000000000_000000100001_100001000001_001010110110_111000000000",	-- 1247
        b"010010001000_000000000000_000000100001_110001010100_001010110011_111000000000",	-- 1250
        b"100101101000_010000000000_010010100001_110001010111_001010110011_111000000000",	-- 1251
        b"100101101000_010000000000_010010100001_110001010011_001010110011_111000000000",	-- 1252
        b"100101101000_010000000000_010010100001_110001011000_001010110011_111000000000",	-- 1253
        b"110010110000_010001000000_000001101001_111010000010_000000000000_111000000000",	-- 1254
        b"010001101001_010000100000_000000100001_110011000001_001011000110_111000000000",	-- 1255
        b"110010000000_000000000001_011000100001_101010000001_000000000000_111000000000",	-- 1256
        b"110010000000_000000000001_111000100001_101010000001_000000000000_111000000000",	-- 1257
        b"110010000000_000000000001_101000100001_101010000001_000000000000_111000000000",	-- 1260
        b"110010000000_000000000001_001000100001_101010000001_000000000000_111000000000",	-- 1261
        b"110010000000_000000000000_011000100001_101010000001_000000000000_111000000000",	-- 1262
        b"010001101000_010000000010_000000100001_111010000001_000000000000_111000000000",	-- 1263
        b"010010001000_000000000000_000110100001_101110000000_001111111111_111000100000",	-- 1264
        b"011001101000_010000000000_000000100001_101010000001_000000000000_111000000000",	-- 1265
        b"010010000000_000000000000_000000100001_001110000000_000000000000_111010000000",	-- 1266
        b"110010110000_010000100000_000001101001_111010000010_000000000000_111000000000",	-- 1267
        b"110010000000_000000000000_000000100001_100011000001_001011000110_111000000000",	-- 1270
        b"010010001000_000000000000_000000100001_101110000000_001011000001_111000100000",	-- 1271
        b"010010001000_000100100000_000000100001_110001000001_101000001110_111000000000",	-- 1272
        b"010001101111_111011011000_000000100001_111110000000_000000000000_111000000000",	-- 1273
        b"110010000000_000000000000_000110100001_101110000000_000100100101_111000100000",	-- 1274
        b"010001101011_011011011010_000000100001_110001000001_100111000100_111010000000",	-- 1275
        b"010001101011_011011011000_001010100001_110001000001_100101111011_001001000000",	-- 1276
        b"110001101100_110000000000_000001101001_110011000010_001010111100_111000000000",	-- 1277
        b"110010000000_000000000000_000000100001_100011000001_000100111111_111000000000",	-- 1300
        b"011011000111_110000000000_000000100001_101110000000_000000000000_111000000000",	-- 1301
        b"110010111101_111000000000_000001101001_110011000010_000101001001_111000000000",	-- 1302
        b"110010000000_000000000000_000000100001_100011000001_000100111111_111000000000",	-- 1303
        b"010010001000_000000000000_000000100001_101110000000_001000000000_111000100000",	-- 1304
        b"110010000000_000000000000_000000100001_101011000001_001001110110_111000000000",	-- 1305
        b"011001101110_010000000000_000000100001_101110000000_000000000000_111000000000",	-- 1306
        b"110001101000_010000100000_000000100001_110011000001_001011000111_111000000000",	-- 1307
        b"110001101110_110000000001_110100100001_111101000001_000000000000_111000000000",	-- 1310
        b"010011000110_111011100000_000000100001_111101000001_000000000000_111000000000",	-- 1311
        b"110010000000_000000000000_000110100001_101101000001_000101101101_111000100000",	-- 1312
        b"110011000111_111011011000_000000100001_111101000001_000000000000_111010000000",	-- 1313
        b"110010000000_000000000000_000110100001_101110000000_000101101011_111000100000",	-- 1314
        b"010010000000_000011011000_000001101001_100011000010_001100000001_111010000000",	-- 1315
        b"110010000000_000000000000_000110100001_101110000000_000101101100_111000100000",	-- 1316
        b"010010001000_000000000000_000000100001_101110000000_001100001101_111000100000",	-- 1317
        b"110011000111_111100100000_000000100001_110001000001_101000010001_111010000000",	-- 1320
        b"010010001000_000000000000_000000100001_110001011100_001010110011_111000000000",	-- 1321
        b"100101101000_010000000000_010010100001_110001011110_001010110011_111000000000",	-- 1322
        b"100101101000_010000000000_010010100001_110001100000_001010110011_111000000000",	-- 1323
        b"100101101000_010000000000_010010100001_110001100010_001010110011_111000000000",	-- 1324
        b"100101101000_010000000000_010010100001_110001100100_001010110011_111000000000",	-- 1325
        b"100101101000_010000000000_010010100001_110001100110_001010110011_111000000000",	-- 1326
        b"100101101000_010000000000_010010100001_110001110110_001010110011_111000000000",	-- 1327
        b"010001101000_010100100000_000000100001_110001000001_100111000100_111000000000",	-- 1330
        b"010001101000_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1331
        b"010001101001_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1332
        b"010001101001_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1333
        b"010001101010_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1334
        b"010001101010_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1335
        b"010001101011_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1336
        b"010001101011_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1337
        b"010001101100_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1340
        b"110010000000_000000000000_000110100001_101110000000_000101101100_111000100000",	-- 1341
        b"010010000000_000100100000_000000100001_100001000001_100111000011_111010000000",	-- 1342
        b"010001101101_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1343
        b"010001101101_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1344
        b"010001101110_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1345
        b"010001101110_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1346
        b"010001101111_010100100000_000000100001_110001000001_100111000011_111000000000",	-- 1347
        b"010001101111_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1350
        b"010001101000_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1351
        b"010001101000_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1352
        b"010001101001_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1353
        b"010001101001_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1354
        b"010001101010_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1355
        b"010001101010_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1356
        b"110010000000_000000000000_000110100001_101110000000_000101101101_111000100000",	-- 1357
        b"010010000000_000100100000_000000100001_100001000001_100111000011_111010000000",	-- 1360
        b"010001101011_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1361
        b"010001101100_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1362
        b"010001101100_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1363
        b"010001101101_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1364
        b"010001101101_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1365
        b"010001101110_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1366
        b"010001101110_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1367
        b"010001101111_011100100000_000000100001_110001000001_100111000011_111000000000",	-- 1370
        b"010001101111_111100100000_000000100001_110001000001_100111000011_111000000000",	-- 1371
        b"010010001000_000010000000_000110100001_101110000000_000001101001_111000100000",	-- 1372
        b"010010001000_000010100000_000000100001_101110000000_000000001001_111000100000",	-- 1373
        b"010010000000_000100100000_000000100001_100001000001_100111000011_111010000000",	-- 1374
        b"010001101010_010010000010_000110100001_111110000000_000000000000_111000000000",	-- 1375
        b"010010000000_000100100000_000000100001_101110000000_000000000000_111010000000",	-- 1376
        b"110010001000_000000000000_000000100001_110001000001_100111000011_111010000000",	-- 1377
        b"010000110111_111010100000_000001101001_110011000011_001011111101_111000000000",	-- 1400
        b"010010001000_000000000000_000000100001_110001000001_001010100000_111000000000",	-- 1401
        b"010001101100_111000000000_011000100001_101110000000_000000000011_111000100000",	-- 1402
        b"110010000000_000000000000_000000100001_100001000001_000111100011_111000000000",	-- 1403
        b"010010001000_000010100000_000000100001_101110000000_000001001000_111000100000",	-- 1404
        b"110010000000_000000000000_000000100001_100001000001_000101101110_111000000000",	-- 1405
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 1406
        b"010010000000_000000000000_000000100001_100001000001_000101011011_111010000000",	-- 1407
        b"110010000000_000000000000_000000100001_100001000001_000101110101_111000000000",	-- 1410
        b"010001101000_011000000000_000000100001_110001000001_000101100000_111000000000",	-- 1411
        b"110010000000_000000000000_000000100001_100001000001_000101110101_111000000000",	-- 1412
        b"010001101011_110000000000_000000100001_110001000001_000101011011_111000000000",	-- 1413
        b"110010000000_000000000000_000000100001_100011000001_000011100001_111000000000",	-- 1414
        b"010010001000_000000000000_000000100001_101110000000_000000000101_111000100000",	-- 1415
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 1416
        b"110011000111_111000000000_000000100001_110011000001_001100000001_111010000000",	-- 1417
        b"110010000000_000000000000_000000100001_100011011101_001011000100_111000000000",	-- 1420
        b"110010000000_000000000000_000000100001_100001000001_000011101110_111000000000",	-- 1421
        b"011101101011_110100000001_111110100001_111011100011_001011001000_111000000000",	-- 1422
        b"011011001111_010000000001_100000100001_001011111010_001100010111_111010000000",	-- 1423
        b"010011111000_010011011000_001010100001_111011011000_001100011001_001001000000",	-- 1424
        b"010001101011_110011110010_000000100001_110001000001_100110110010_111000000000",	-- 1425
        b"110010000000_000000000000_000000100001_101011000001_001100011101_111000000000",	-- 1426
        b"010001101100_010011011000_100110100001_111011010011_001100010101_111000000000",	-- 1427
        b"010001101100_010011011000_001010100001_111110000000_000000000000_001001000000",	-- 1430
        b"010001101011_110011110010_000000100001_110001010001_100001101100_000000000000",	-- 1431
        b"010010000000_000011000000_110110100001_001110000000_000000000000_101100100000",	-- 1432
        b"010001101011_010100010000_000000100001_111011110001_001100011110_000000000000",	-- 1433
        b"010000110111_111011110000_000000100001_110011000001_001100010101_111000000000",	-- 1434
        b"010001101100_110011000000_110110100001_111110000000_000000000000_111100100000",	-- 1435
        b"010001101011_010100010000_101110100001_110110001010_100000000000_111000000000",	-- 1436
        b"110001101011_010000000000_110110100001_110001000001_001100101000_111000000000",	-- 1437
        b"110010000000_000000000000_101110100001_100110000001_100000000000_111000000000",	-- 1440
        b"010010001000_000110010000_000000100001_101110000000_000100000000_111000100000",	-- 1441
        b"010011000110_111100000000_011000100001_110001000001_010100011010_111000000000",	-- 1442
        b"010001101011_010100010000_110110100001_111110000000_000000000000_111000000000",	-- 1443
        b"110010000000_000000000000_000000100001_100001001011_001100101000_111000000000",	-- 1444
        b"110010000000_000000000000_000000100001_100001000001_010100010100_111000000000",	-- 1445
        b"110010000000_000000000000_101110100001_100110000001_100000000000_111000000000",	-- 1446
        b"010001101100_110100010000_011000100001_111010001010_000000000000_111000000000",	-- 1447
        b"011101101111_011000000000_000000100001_100011000100_001100110010_111010000000",	-- 1450
        b"010010000000_000100100000_000000100001_101110000000_000000000000_111010000000",	-- 1451
        b"110011001000_010000000000_000000100001_010011010111_001100110001_111000000000",	-- 1452
        b"011010010111_110100000000_000001000001_100011000010_001100110001_111000000000",	-- 1453
        b"010000111000_010100000000_010000100001_110011101111_001100101111_111000000000",	-- 1454
        b"010000110111_110100000000_000000100001_111010001001_000000000000_111000000000",	-- 1455
        b"110010000000_000000000000_000000100001_100011000001_001100110010_111000000000",	-- 1456
        b"110010000000_000000000000_000000100001_101010001001_000000000000_111000000000",	-- 1457
        b"110010000000_000000000000_000000100001_100011000001_001100110010_111000000000",	-- 1460
        b"010000110000_010100010000_011000100001_111010001001_000000000000_111000000000",	-- 1461
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 1462
        b"010010000000_000000000000_000000100001_100011010111_001100100111_111010000000",	-- 1463
        b"110010000000_000000000000_010000100001_101011001100_100111100111_111000000000",	-- 1464
        b"110010000000_000000000000_000000100001_100011001111_001100100111_111000000000",	-- 1465
        b"010001101100_110100000001_111110100001_111010001010_000000000000_111000000000",	-- 1466
        b"011000110100_110000000000_000000100001_100011000100_001100110010_111000000000",	-- 1467
        b"010011001111_111100000001_111110100001_111010001001_000000000000_111000000000",	-- 1470
        b"110010000000_000000000000_000000100001_100011000001_001100110010_111000000000",	-- 1471
        b"010010000000_000101100000_101110100001_001110000000_000000010000_111010000000",	-- 1472
        b"010010000000_000001011000_101110100001_100110000001_100100000000_111010000000",	-- 1473
        b"010010000000_000101000000_101110100001_101110000000_000000010000_111010000000",	-- 1474
        b"010010000000_000000111000_000000100001_100011000001_001100111110_111010000000",	-- 1475
        b"011111000110_111100000001_111110100001_110011100110_001101000010_111000000000",	-- 1476
        b"110010000000_000000000000_000000100001_100001000001_100110110011_111000000000",	-- 1477
        b"010001101100_110101100000_000000100001_110001000001_100110110000_111000000000",	-- 1500
        b"010001101100_110001011000_000000100001_110011000001_001101000111_111000000000",	-- 1501
        b"010010001000_000110010000_000000100001_101110000000_000010000000_111000100000",	-- 1502
        b"110010000000_000000000000_000000100001_100001000001_010100011010_111000000000",	-- 1503
        b"011111000110_111100000001_111110100001_110001000001_100110110011_111000000000",	-- 1504
        b"010001101100_110101100000_000000100001_110001000001_100110110000_111000000000",	-- 1505
        b"010001101100_110001011000_000000100001_110001000001_010100010100_111000000000",	-- 1506
        b"110001101101_110000000000_101110100001_010110000001_100100000000_111000000000",	-- 1507
        b"010010000000_000101000000_000000100001_100011000001_001101001001_111010000000",	-- 1510
        b"011101101100_010011011001_111110100001_110001100111_100110110011_111000000000",	-- 1511
        b"011101101100_110101100000_101110100001_010110100111_100100000000_111000000000",	-- 1512
        b"110010000000_000000000000_000000100001_100001000001_010100010001_111000000000",	-- 1513
        b"011101101100_110101100000_101110100001_010110000001_100100000000_111000000000",	-- 1514
        b"010010000000_000101000000_000000100001_100011000001_001101001110_111010000000",	-- 1515
        b"011101101100_010100000001_111110100001_110001100111_100110110011_111000000000",	-- 1516
        b"011101101100_110101100000_000000100001_010011100111_001101010010_111000000000",	-- 1517
        b"110010000000_000000000000_000000100001_100001000001_010100010001_111000000000",	-- 1520
        b"011101101100_110101100000_101110100001_011110000000_000000000000_111000000000",	-- 1521
        b"110010000000_000000000000_101110100001_100110101000_100100000000_111000000000",	-- 1522
        b"110010000000_000000000000_000000100001_100110111010_100100000000_111000000000",	-- 1523
        b"110010000000_000000000000_000000100001_100001000001_100111011000_111000000000",	-- 1524
        b"110010000000_000000000000_101110100001_100110000001_100100000000_111000000000",	-- 1525
        b"010010000000_000101000000_000000100001_100011000001_001101010111_111010000000",	-- 1526
        b"010010000111_110101100000_000000100001_101110000000_000000000000_111011100000",	-- 1527
        b"011111000100_010101100000_101110100001_010110000001_100100000000_111000000000",	-- 1530
        b"010010000000_000101100000_000000100001_100110000001_100100000000_111010000000",	-- 1531
        b"010010000000_000101100000_000000100001_101110000000_000000000000_111010000000",	-- 1532
        b"010001101101_110101100000_000000100001_010110000001_100100000000_111000000000",	-- 1533
        b"010010000000_000101000000_000000100001_101110000000_000000000000_111010000000",	-- 1534
        b"110010000000_000000000000_000000100001_100001000001_001101100000_111000000000",	-- 1535
        b"110010000000_000000000000_101110101101_100110000011_101000000000_111000000000",	-- 1536
        b"110010000000_000000000000_000000100001_100011000001_100111100101_111000000000",	-- 1537
        b"010011000110_111100000000_000000011110_110001000001_001101100101_111000000000",	-- 1540
        b"010001101100_010011011000_001011011101_110011000010_001101110010_011001000000",	-- 1541
        b"010010000000_000101100000_000000100001_001110000000_000000000000_101001000000",	-- 1542
        b"110010000000_000000000000_000000011100_101010110001_000000000000_111000000000",	-- 1543
        b"110010000000_000000000000_000000011110_101010000001_000000000000_111000000000",	-- 1544
        b"010010001000_000000000000_000000100001_101110000000_111111110000_111000100000",	-- 1545
        b"010010000000_010000000000_000000011110_101110000000_000000000000_111011100000",	-- 1546
        b"110011000000_010100000000_000001101001_111011000011_001101101001_111000000000",	-- 1547
        b"010010001000_000000000000_000000100001_101110000000_000011000000_111000100000",	-- 1550
        b"110000100100_010000000000_000001111101_011010000011_000000000000_111000000000",	-- 1551
        b"010001101100_010010100000_000110100001_111110000000_000000000000_111000000000",	-- 1552
        b"000101101010_110001000000_000010100001_110100000001_000000000001_111000000000",	-- 1553
        b"000101101001_010001000000_000010100001_111000000000_000000000000_111000000000",	-- 1554
        b"010010001000_000000100000_000000100001_101110000000_000000000111_111000100000",	-- 1555
        b"010010010000_110010100000_000000100001_111110000000_000000000000_111000000000",	-- 1556
        b"010011000000_110001000000_000000100001_111110000000_000000000000_111000000000",	-- 1557
        b"010010000001_010010101000_000000100001_101110000000_000000000000_111011100000",	-- 1560
        b"010010001000_000000000000_000000100001_101010000001_000001111111_111000100000",	-- 1561
        b"011000100100_010000000010_000001111101_011010000010_000000000000_111000000000",	-- 1562
        b"010010000000_000101100000_000001001001_100011000010_001101111111_111010000000",	-- 1563
        b"110010000000_000000000000_000000011100_101110000000_000000000000_111000000000",	-- 1564
        b"011011000000_110010100000_000001101001_111010000011_000000000000_111000000000",	-- 1565
        b"110010000000_000000000000_000000100001_100001000001_011111000111_111000000000",	-- 1566
        b"010010001000_000000100000_000000100001_101110000000_000011000000_111000100000",	-- 1567
        b"010011000000_110000000000_000000100001_110001000001_100000010111_111000000000",	-- 1570
        b"010010010000_110101100000_000000100001_110001000001_100000010110_111000000000",	-- 1571
        b"010011110000_010101100000_000000100001_111010000001_000000000000_111000000000",	-- 1572
        b"010010000000_000101100000_000000011100_100001000001_011100001110_111010000000",	-- 1573
        b"010010010000_010010100000_000110100001_111110000000_000000000000_111000000000",	-- 1574
        b"010010000000_000010000000_000000100001_100001000001_011110110101_111010000000",	-- 1575
        b"110010000000_000000000000_000000100001_100011000001_011010010101_111000000000",	-- 1576
        b"010010000000_000101100000_000000011100_101010000001_000000000000_111010000000",	-- 1577
        b"110010000000_000000000000_000000100001_100011010111_001110001010_111000000000",	-- 1600
        b"110010000000_000000000000_000000100001_100011011111_001110011111_111000000000",	-- 1601
        b"010010001000_000011011000_000000100001_101110000000_000100010000_111000100000",	-- 1602
        b"010000110010_011011011000_001010100001_110001000001_100101111011_001001000000",	-- 1603
        b"010001101100_110011011000_010000100001_110001000001_001110010101_111000000000",	-- 1604
        b"011101101011_011100000001_111110100001_110001000001_100111001010_111000000000",	-- 1605
        b"010001101011_110100100000_000000100001_110001000001_100111001000_111000000000",	-- 1606
        b"010001101101_110100100000_000000100001_110001000001_100111001000_111000000000",	-- 1607
        b"010001101100_010100000011_111110100001_110001000001_100110110011_111000000000",	-- 1610
        b"010001101100_110011100000_011000100001_111011000001_001100010000_111000000000",	-- 1611
        b"010010000011_010100100000_000000100001_100001000001_001110011101_111011100000",	-- 1612
        b"010010000100_010100101000_000000100001_100001000001_001110010100_111011100000",	-- 1613
        b"010010001000_000100000000_000000100001_101110000000_000000100000_111000100000",	-- 1614
        b"010001101100_010011011000_000000100001_110011011111_001110010001_111000000000",	-- 1615
        b"011101101100_010100000001_111110100001_110001000001_100111001010_111000000000",	-- 1616
        b"011101101100_010100000011_111110100001_110001000001_100110110011_111000000000",	-- 1617
        b"110010000000_000000000000_000000100001_101011000001_001100011101_111000000000",	-- 1620
        b"010000110001_111011011000_000000100001_110001000001_100111000100_111000000000",	-- 1621
        b"010001101011_011011011010_001010100001_110001000001_100101111011_001001000000",	-- 1622
        b"110010000000_000000000000_000000100001_100011000001_001100011101_111000000000",	-- 1623
        b"010010000100_110100100000_000000100001_101010000001_000000000000_111011100000",	-- 1624
        b"010010000011_010100100000_000000100001_100001000001_001110011101_111011100000",	-- 1625
        b"010001101000_011100101000_000000100001_111110000000_000000000000_111000000000",	-- 1626
        b"010011000110_111011100000_000000100001_111110000000_000000000000_111000000000",	-- 1627
        b"010001101100_010101100001_111110100001_111110000000_000000000000_111000000000",	-- 1630
        b"010011000110_111101100000_000000100001_111010010010_000000000000_111000000000",	-- 1631
        b"110001101011_110000000001_111110100001_111010011101_000000000000_111000000000",	-- 1632
        b"110010000000_000000000000_000000100001_101010010111_000000000000_111000000000",	-- 1633
        b"010001101101_111101101000_000000100001_111010000001_000000000000_111000000000",	-- 1634
        b"010010001000_000000000000_000000100001_101110000000_000000011111_111000100000",	-- 1635
        b"010010010000_010100100000_000000100001_111010000001_000000000000_111000000000",	-- 1636
        b"010010001000_000011011000_000000100001_101101000001_000100010100_111000100000",	-- 1637
        b"010000110010_011011011000_000000100001_110001000001_001110010101_111000000000",	-- 1640
        b"110010000000_000000000000_000000100001_100011100100_001110101001_111000000000",	-- 1641
        b"010010000100_110100100000_000000100001_101110000000_000000000000_111011100000",	-- 1642
        b"010001101100_010100110000_000000100001_110001000001_100111000100_111000000000",	-- 1643
        b"010001101000_011100100000_000000100001_111110000000_000000000000_111000000000",	-- 1644
        b"010001101011_110100110000_000000100001_110001000001_100111000011_111000000000",	-- 1645
        b"110010000000_000000000000_000000100001_100001000001_011011110000_111000000000",	-- 1646
        b"110010000000_000000000000_000000100001_100001000001_100111000011_111000000000",	-- 1647
        b"010001101011_011011011010_000000100001_110011000001_001110101110_111000000000",	-- 1650
        b"010011000110_111011100000_000000100001_110001000001_100111000100_111000000000",	-- 1651
        b"010001101011_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1652
        b"010001101101_110100100000_000000100001_110001000001_100111000011_111000000000",	-- 1653
        b"110010000000_000000000000_000000100001_100001000001_011011110000_111000000000",	-- 1654
        b"011101101011_011011011000_000000100001_110001000001_100111000011_111000000000",	-- 1655
        b"010010001000_000000011000_000000100001_110011011111_001110110011_111000000000",	-- 1656
        b"010010001000_000000000000_100000100001_101101000001_000000000100_111000100000",	-- 1657
        b"010000110000_010011011000_000000100001_111101000001_000000000000_111000000000",	-- 1660
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 1661
        b"010010000000_010000011000_000000100001_101110000000_000000000000_111011100000",	-- 1662
        b"010001101011_011011011010_001010100001_110001000001_100101111011_001001000000",	-- 1663
        b"010001101100_110011100000_011000100001_110011100100_001100010000_111000000000",	-- 1664
        b"010011110000_011100100000_000000100001_110011000001_010011001101_111000000000",	-- 1665
        b"011000110001_011001011000_000000100001_101110000000_000000000000_111000000000",	-- 1666
        b"011001011000_000000000010_000000100001_011110000000_000000000000_111000000000",	-- 1667
        b"010001111101_110101100000_000001010100_111110000000_000000000000_111000000000",	-- 1670
        b"000111001111_111001011000_000011001001_110110000011_101000000000_111000000000",	-- 1671
        b"110010000000_000000000000_000000101001_100011000010_010000111101_111000000000",	-- 1672
        b"110010000000_000000000000_000000101101_100110000011_101000000000_111000000000",	-- 1673
        b"110010000000_000000000000_000000100001_100011000001_010000111000_111000000000",	-- 1674
        b"010001101101_010000111000_000000100001_010011000110_100001010111_111000000000",	-- 1675
        b"110001101010_110000000000_000001011101_010011000010_001111000000_111000000000",	-- 1676
        b"010010001000_000101000000_000000100001_110011000001_001111000001_111000000000",	-- 1677
        b"010000001000_000101000000_000000100001_111110000000_000000000000_111000000000",	-- 1700
        b"011010010111_110010000000_000001001001_000011000010_001111010111_111000000000",	-- 1701
        b"011000011010_110000000010_000001111101_100011000011_001111000010_111000000000",	-- 1702
        b"010010001000_000000000000_000000100001_101110000000_000000100100_111000100000",	-- 1703
        b"010000001000_000001000000_000000100001_011110000000_000000000000_111000000000",	-- 1704
        b"011000111010_110000000000_000000100001_101110000000_000000000000_111000000000",	-- 1705
        b"110000101000_010000000010_000001111101_110011000010_001111001000_111000000000",	-- 1706
        b"010001101001_010001000010_000000100001_010011000001_001111000101_111000000000",	-- 1707
        b"010001101101_010000111000_000001000001_010011000010_010001101111_111000000000",	-- 1710
        b"010001101001_010101100000_000000100001_010001000001_010001010110_111000000000",	-- 1711
        b"110001101001_011000000000_000001101000_110011000010_001111001011_111000000000",	-- 1712
        b"000101101010_010101000001_010010100001_110100000001_000000000100_111000000000",	-- 1713
        b"000101101101_010101000001_010010100001_111000000000_000000000000_111000000000",	-- 1714
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 1715
        b"010010000000_010000000000_101110100001_101110000000_000000000000_111011100000",	-- 1716
        b"110011000000_010101000000_000001101001_100011000011_001111010001_111000000000",	-- 1717
        b"010000110101_110101010000_000000100001_111011000001_100011101000_111000000000",	-- 1720
        b"110010000000_000000000000_000000100001_100001000001_100110110000_111000000000",	-- 1721
        b"010000110100_110101100000_101110100001_111110000000_000000010000_111000000000",	-- 1722
        b"010011000110_111101100000_000000100001_111110000000_000000000000_111000000000",	-- 1723
        b"010010010110_111100100000_000000100001_111110000000_000000000000_111000000000",	-- 1724
        b"110011110101_110100100000_101110100001_111110000000_000000000000_111010000000",	-- 1725
        b"110011000111_111101000000_011000100001_111011000001_001100010000_111010000000",	-- 1726
        b"110010000000_000000000000_101110101001_100110000011_101100010000_111000000000",	-- 1727
        b"110011000111_111001011000_000000100001_110110000001_101100000000_111010000000",	-- 1730
        b"110010000000_000000000000_000000100001_100011000110_001111110001_111000000000",	-- 1731
        b"100101101101_110010000000_010010100001_111100000000_000000000001_111000000000",	-- 1732
        b"100100110010_010010000000_010010100001_111001000000_001111011011_111000000000",	-- 1733
        b"011000110010_010010000000_000000100001_101110000000_000000000000_111000000000",	-- 1734
        b"101101101101_110010000001_010010100001_111100000000_000000000100_111000000000",	-- 1735
        b"101101101010_010010000001_010010100001_111001000000_001111011110_111000000000",	-- 1736
        b"010011000110_110010000000_000000100001_111110000000_000000000000_111000000000",	-- 1737
        b"011111001110_110010100000_000000100001_110011010111_001111100100_111000000000",	-- 1740
        b"110011000101_011101100000_000001101001_110011000010_001111100100_111000000000",	-- 1741
        b"011101101100_010100010010_000000010010_110011011100_001111100101_111000000000",	-- 1742
        b"010011001111_111100000000_000000100001_110011000001_001111100101_111000000000",	-- 1743
        b"110001101101_110000000000_110110010000_111100000000_001100100111_111000000000",	-- 1744
        b"110010000000_000000000000_000000101001_100101000010_001100110010_111000000000",	-- 1745
        b"110010000000_000000000000_000000100001_100011100111_001111101010_111000000000",	-- 1746
        b"010010001000_000110010000_000000100001_101110000000_000001000000_111000100000",	-- 1747
        b"110010000000_000000000000_000000100001_100001000001_010100010010_111000000000",	-- 1750
        b"110010000000_000000000000_000000100001_100011000001_001111101011_111000000000",	-- 1751
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 1752
        b"010010001000_000000000000_000000100001_101110000000_000000000000_111000100000",	-- 1753
        b"110000110000_010010100000_000110100001_111110000000_000000000000_111000000000",	-- 1754
        b"110000110111_111010000000_000000100001_011110000000_000000000000_111000100000",	-- 1755
        b"010010000000_000000100000_101110100001_101110000000_000000000000_111010000000",	-- 1756
        b"110010000000_000000000000_000000100001_100110000001_101100000000_111000000000",	-- 1757
        b"110011000100_111000011000_000001101001_110011000011_001111011010_111000000000",	-- 1760
        b"100101101101_110010000000_010010100001_111100000000_000000000001_111000000000",	-- 1761
        b"100100110010_010010000000_010010100001_111001000000_001111110010_111000000000",	-- 1762
        b"011000110010_010010000000_000000100001_101110000000_000000000000_111000000000",	-- 1763
        b"011110011110_111010100000_000000100001_111110000000_000000000000_111000000000",	-- 1764
        b"010000101101_110101100010_000001110101_110011000010_010000000110_111000000000",	-- 1765
        b"000110001000_000000000000_001010100001_101110000000_000000000100_111000100000",	-- 1766
        b"010011000110_111101100000_000000100001_110100000001_000000000010_111000000000",	-- 1767
        b"000101101000_010000000001_010010100001_111000000000_000000000000_111000000000",	-- 1770
        b"010011110000_010101100000_000000100001_111110000000_000000000000_111000000000",	-- 1771
        b"010000101101_110101100010_000000100001_110011010111_010000000101_111000000000",	-- 1772
        b"110011000101_011101100000_000001101001_110011000010_010000000101_111000000000",	-- 1773
        b"011101101100_010100010010_000000100001_110011011100_001111111110_111000000000",	-- 1774
        b"010011001111_111100000000_000000100001_111110000000_000000000000_111000000000",	-- 1775
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 1776
        b"011010010110_111100100000_000000100001_101110000000_000000000000_111000000000",	-- 1777
        b"010001101100_110100100010_000000100001_111110000000_000000000000_111000000000",	-- 2000
        b"010011000110_111100100000_000000100001_111110000000_000000000000_111000000000",	-- 2001
        b"010011111100_110100100000_000000100001_110001000001_100111001001_111000000000",	-- 2002
        b"011100110111_111100010000_000000100001_110011011100_010000000110_111000000000",	-- 2003
        b"010011001111_111100000000_000000100001_110011000001_010000000110_111000000000",	-- 2004
        b"010001101101_110101110010_000000100001_111110000000_000000000000_111000000000",	-- 2005
        b"010001101101_110100100000_000000100001_110001000001_100111001001_111000000000",	-- 2006
        b"011001101010_110000000000_000000100001_100110000001_101000000000_111000000000",	-- 2007
        b"010011110100_111000011000_000000100001_110011000001_001111011101_111000000000",	-- 2010
        b"110010000000_000000000000_000001011101_100011000010_010000010000_111000000000",	-- 2011
        b"010010001000_000000000000_000000100001_101110000000_000000010010_111000100000",	-- 2012
        b"110000100010_010000000000_000001111101_010011000010_010000001111_111000000000",	-- 2013
        b"010010000100_110100100000_000000100001_101110000000_000000000000_111011100000",	-- 2014
        b"010010001000_000100101000_000001001001_110011000010_010000010000_111000000000",	-- 2015
        b"110000100010_010000000000_000000100001_111110000000_000000000000_111000100000",	-- 2016
        b"000101101100_110100100000_000010100001_111001000000_010000001111_111000000000",	-- 2017
        b"110011000100_110000100000_000000100001_111011000001_010000011111_111010000000",	-- 2020
        b"010011000000_110101000000_000001011101_110011000010_010000011011_111000000000",	-- 2021
        b"010010001000_000000000000_000000100001_101110000000_000000010010_111000100000",	-- 2022
        b"110000100010_010000000000_000001111101_010011000010_010000011000_111000000000",	-- 2023
        b"010010000101_010101000000_000000100001_101110000000_000000000000_111011100000",	-- 2024
        b"010010001000_000101010000_000000100001_110001000001_100000010111_111000000000",	-- 2025
        b"010010001000_000000110000_000001001001_110011000010_010000011000_111000000000",	-- 2026
        b"110000100010_010000000000_000000100001_111110000000_000000000000_111000100000",	-- 2027
        b"011001101000_110000000000_000000100001_101110000000_000000000000_111000000000",	-- 2030
        b"101101101101_010101000000_010010100001_111001000000_010000011001_111000000000",	-- 2031
        b"010011001111_111000100000_000000100001_111110000000_000000000000_111000000000",	-- 2032
        b"010010010000_110100100000_000000100001_110011100111_010000011110_111000000000",	-- 2033
        b"010011110101_010100100000_000000100001_110001000001_010100001100_111000000000",	-- 2034
        b"110010000000_000000000000_000000100001_100011000001_010000011111_111000000000",	-- 2035
        b"010011110101_010100100000_000000100001_110001000001_100111001001_111000000000",	-- 2036
        b"010010010100_111000011000_011000100001_111011000001_001100010000_111000000000",	-- 2037
        b"100101101101_110101100000_010011011101_110011000011_010000100010_111000000000",	-- 2040
        b"010001111101_110101100010_000000100001_111110000000_000000000000_111000000000",	-- 2041
        b"100101101101_110101100001_010010100001_110100000001_000000000110_111000000000",	-- 2042
        b"100101101101_110101100001_010010100001_111000000000_000000000000_111000000000",	-- 2043
        b"011011000111_010101100000_011000100001_101110000000_000000000000_111000000000",	-- 2044
        b"010010010111_010101100000_000000100001_111110000000_000000000000_111000000000",	-- 2045
        b"010010001000_000000100000_000000100001_101110000000_000010100010_111000100000",	-- 2046
        b"110000101000_110000000010_000000100000_111110000000_000000000000_111000100000",	-- 2047
        b"110010000000_000000000000_000000111101_100011000010_010001110001_111000000000",	-- 2050
        b"001111000111_111101100000_110010101001_110011000010_010000101011_111000000000",	-- 2051
        b"001111000111_111101100000_110010100001_111001000000_010000101010_111000000000",	-- 2052
        b"110011000111_111101100000_000001011101_110110000011_101000000000_111010000000",	-- 2053
        b"010001111101_110101100010_000000100001_110110000001_101000000000_111010000000",	-- 2054
        b"110011001111_111000000000_000001111101_111011000011_001100010000_111000000000",	-- 2055
        b"110001101101_110000000010_000001011101_111011000011_001100010000_111010000000",	-- 2056
        b"110000110111_111101100000_000000100001_111011000001_001100010000_111010000000",	-- 2057
        b"110010000000_000000000000_000000100001_100011000001_100011100011_111000000000",	-- 2060
        b"110010010111_110100000000_011000100001_111011000001_001100010000_111010000000",	-- 2061
        b"010010000100_010100000000_101110100001_101110000000_000000000000_111011100000",	-- 2062
        b"110011000111_110100000000_011000100001_110011000001_001100010000_111010000000",	-- 2063
        b"010010000101_110101100000_000000100001_100110000001_101000000000_111011100000",	-- 2064
        b"110010000000_000000000000_000001011101_100110000011_101000000000_111000000000",	-- 2065
        b"010001111101_110101100010_000001101000_110011000010_010000111101_111000000000",	-- 2066
        b"110010000000_000000000000_000001001101_100110000011_101000000000_111000000000",	-- 2067
        b"010010001000_000000000001_111000100001_101110000000_101000000010_111000100000",	-- 2070
        b"010010000000_010000000000_000000100001_100001000001_100001101001_111011100000",	-- 2071
        b"110010000000_000000000000_101110100001_100110000001_101000000000_111000000000",	-- 2072
        b"010000110101_010101100000_000001101101_010011000010_010000111111_111000000000",	-- 2073
        b"110010000000_000000000000_000001010111_100110000010_101000000000_111000000000",	-- 2074
        b"010011110110_011000011000_101110100001_110110000001_101000000000_111000000000",	-- 2075
        b"010000100101_010101100000_000001101111_010011000010_010000111100_111000000000",	-- 2076
        b"110010000000_000000000000_000001010111_100011000010_010000111000_111000000000",	-- 2077
        b"010010001000_000000000001_111000100001_101110000000_110000000010_111000100000",	-- 2100
        b"010010000000_010000000000_000000100001_100001000001_100001101001_111011100000",	-- 2101
        b"110010000000_000000000000_101110100001_100110000001_101000000000_111000000000",	-- 2102
        b"010010001000_000101100000_000000100001_111100000000_000000100001_111000000000",	-- 2103
        b"001000000101_010101100000_110010100001_111110000000_000000000000_111000000000",	-- 2104
        b"001000000101_010101100000_110010100001_111001000000_010001000101_111000000000",	-- 2105
        b"011000000101_010101100100_110010100001_111110000000_000000000000_111000000000",	-- 2106
        b"101001101101_110101100000_100010100001_011110000000_000000000000_111000000000",	-- 2107
        b"000111001111_111001011000_101011011101_110110000010_101000000000_111000000000",	-- 2110
        b"110010000000_000000000000_000001010101_100110000011_101000000000_111000000000",	-- 2111
        b"000110001000_000101100000_001010100001_110001000001_100001100011_111000000000",	-- 2112
        b"000110001000_000001011000_001010100001_110110000001_101000000000_111000000000",	-- 2113
        b"010001101101_110101100010_000001001001_010011000010_010001001110_111000000000",	-- 2114
        b"110010000000_000000000000_000001001001_100001000011_100001100011_111000000000",	-- 2115
        b"010001101001_011101100000_000000100001_110110000001_101100000000_111000000000",	-- 2116
        b"010001101101_010000111000_000001111101_110011000010_010001010001_111000000000",	-- 2117
        b"010010001000_000101000000_000000100001_110011000001_010001010100_111000000000",	-- 2120
        b"010000001000_000101000000_000000100001_110011000001_010001010100_111000000000",	-- 2121
        b"110010000000_000000000000_101110100001_101110000000_000000010000_111000000000",	-- 2122
        b"010010000000_000000111000_000000100001_101110000000_000000000000_111010000000",	-- 2123
        b"010001101101_110001000000_000000100001_010001000001_010001010110_111000000000",	-- 2124
        b"110010000000_000000000000_000000100001_100110000001_101000000000_111000000000",	-- 2125
        b"010001101101_010000100000_000001011101_010011000011_010001011000_111000000000",	-- 2126
        b"010001111001_010001000010_000000100001_111110000000_000000000000_111000000000",	-- 2127
        b"011000110000_111000111000_000001011101_100011000011_010001011011_111000000000",	-- 2130
        b"110001011000_000000000010_000000100000_101110000000_000000000000_111000000000",	-- 2131
        b"010001111000_110000100110_000000000001_111110000000_000000000000_111000000000",	-- 2132
        b"110000100000_110001000010_000001111101_100011000011_010001101111_111000000000",	-- 2133
        b"001001101101_010101000000_101010100001_111110000000_000000000000_111000000000",	-- 2134
        b"101000000101_110101000001_111010100001_111100000000_000000100001_111000000000",	-- 2135
        b"110000000101_110101000101_111010100001_111110000000_000000000000_111000000000",	-- 2136
        b"110000000101_110101000101_111010100001_111001000000_010001011111_111000000000",	-- 2137
        b"111000000101_110101000100_011010100001_111110000000_000000000000_111000000000",	-- 2140
        b"010001101101_010001011000_000001011100_110011000010_010001100110_111000000000",	-- 2141
        b"110001101101_110000000000_000000111101_010011000011_010001101110_111000000000",	-- 2142
        b"110010000000_000000000000_000001011101_100011000010_010001101001_111000000000",	-- 2143
        b"010000110101_110001011000_000000100001_111110000000_000000000000_111000000000",	-- 2144
        b"010000111111_111101100000_000000100001_111010000001_000000000000_111000000000",	-- 2145
        b"110001101101_110000000000_000000101001_010011000010_010001101110_111000000000",	-- 2146
        b"110000110001_011001000000_000000111100_110011000010_010001101011_111000000000",	-- 2147
        b"110010000000_000000000000_000001011101_100011000010_010001100100_111000000000",	-- 2150
        b"010000010101_110001011010_000000100001_111110000000_000000000000_111000000000",	-- 2151
        b"010001101000_000101100010_000000100001_111010000001_000000000000_111000000000",	-- 2152
        b"110010000000_000000000000_000000101001_100011000011_010001101110_111000000000",	-- 2153
        b"110010000000_000000000000_000001011101_100011000010_010001101001_111000000000",	-- 2154
        b"010000110101_110001011000_000000100001_110011000001_010001100101_111000000000",	-- 2155
        b"010011001111_111101100000_000000100001_111010000001_000000000000_111000000000",	-- 2156
        b"010010001000_000000000000_000000100001_101110000000_000000100000_111000100000",	-- 2157
        b"010010000000_010000000000_000000100001_100001000001_100001101011_111011100000",	-- 2160
        b"110010000000_000000000000_011000100001_100001000001_100001100011_111000000000",	-- 2161
        b"110010000000_000000000000_000000100001_101011000001_100001011000_111000000000",	-- 2162
        b"100101101000_111000111000_010010100001_110001000001_010001111001_111000000000",	-- 2163
        b"010000110000_111001011000_000000100001_011110000000_000000000000_111000000000",	-- 2164
        b"010000110101_010101100000_000001010101_011110000000_000000000000_111000000000",	-- 2165
        b"000101101001_011001011000_101011001101_110011000010_010000111111_111000000000",	-- 2166
        b"110010000000_000000000000_000001010111_100110000010_101000000000_111000000000",	-- 2167
        b"010011110110_011000011000_000000100001_110110000001_101000000000_111000000000",	-- 2170
        b"100101101001_011001011000_010010100001_111010000001_000000000000_111000000000",	-- 2171
        b"100101101000_111000111000_010010100001_110001000001_010001111001_111000000000",	-- 2172
        b"010000100000_111001011000_000000100001_011110000000_000000000000_111000000000",	-- 2173
        b"010000100101_010101100000_000001010101_010011000001_010001110110_111000000000",	-- 2174
        b"110010000000_000000000000_000000100001_100110000001_101000000000_111000000000",	-- 2175
        b"110001101101_110000000000_000000100001_001110000000_000000000000_111000000000",	-- 2176
        b"011000110001_011001011000_000000100001_100011000001_010010000001_111000000000",	-- 2177
        b"011001101001_011000000000_000000100001_100011000001_010010000001_111000000000",	-- 2200
        b"010010001000_000000000000_011000100001_101110000000_000011111111_111000100000",	-- 2201
        b"010011000000_010100000000_000000100000_110011101110_010010000110_111000000000",	-- 2202
        b"010000110111_111100000000_000000100001_111110000000_000000000000_111000100000",	-- 2203
        b"110010000000_000000000000_101110101001_100110000011_101000000000_111000000000",	-- 2204
        b"110010000000_000000000000_011000100001_101011000001_001100010000_111000000000",	-- 2205
        b"010000100000_010100000000_000000100001_111110000000_000000000000_111000100000",	-- 2206
        b"110010000000_000000000000_101110100001_100110000001_101100000000_111000000000",	-- 2207
        b"010000110101_110101100000_000000001100_111001000000_010010001000_111000000000",	-- 2210
        b"110011000111_111101100000_011000101101_111011000011_001100010000_111010000000",	-- 2211
        b"010000110101_110101100000_000000100001_110001000001_100001100011_111000000000",	-- 2212
        b"000101000000_000101100000_101010100001_111011000001_100001011000_111010000000",	-- 2213
        b"000101101101_110101100000_101010100001_111001000000_010010001100_111000000000",	-- 2214
        b"110011000111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2215
        b"001001101101_110101100000_101010100001_111110000000_000000000000_111000000000",	-- 2216
        b"101000000101_110101100000_110010001100_111001000000_010010001111_111000000000",	-- 2217
        b"101101101101_110101100000_110010100001_111110000000_000000000000_111000000000",	-- 2220
        b"101101101101_110101100000_110010100001_111110000000_000000000000_111000000000",	-- 2221
        b"001101000000_000101100000_101010100001_111110000000_000000000000_111010000000",	-- 2222
        b"110010000000_000000000000_101110100001_101110000000_000000010000_111000000000",	-- 2223
        b"000111001111_111001011000_101010101101_110011000011_001100010000_111010000000",	-- 2224
        b"110010000000_000000000000_000000100001_101011000001_010001110001_111000000000",	-- 2225
        b"001001101101_110101100000_101010100001_111001000000_010010010110_111000000000",	-- 2226
        b"110001101101_110000000000_101110100001_111110000000_000000010000_111010000000",	-- 2227
        b"000111001111_111001011000_101010100001_111011000001_001100010000_111010000000",	-- 2230
        b"100101101101_110101100000_010010100001_111001000000_010010011001_111000000000",	-- 2231
        b"110011000111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2232
        b"000101101101_110101100000_000010100001_111001000000_010010011011_111000000000",	-- 2233
        b"110011000111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2234
        b"101101101101_110101100000_110010100001_111001000000_010010011101_111000000000",	-- 2235
        b"010011001111_111001011000_000000100001_110011000001_100011100000_111000000000",	-- 2236
        b"001101101101_110101100000_110010100001_111001000000_010010011111_111000000000",	-- 2237
        b"010011001111_111001011000_000000100001_110011000001_100011100000_111000000000",	-- 2240
        b"100101101101_110101100001_010010100001_111001000000_010010100001_111000000000",	-- 2241
        b"110011000111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2242
        b"000101101101_110101100001_010010100001_111001000000_010010100011_111000000000",	-- 2243
        b"110011000111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2244
        b"101101101101_110101100001_111010100001_111001000000_010010100101_111000000000",	-- 2245
        b"010011001111_111001011000_000000100001_110011000001_100011100000_111000000000",	-- 2246
        b"001101101101_110101100001_111010100001_111001000000_010010100111_111000000000",	-- 2247
        b"010011001111_111001011000_000000100001_110011000001_100011100000_111000000000",	-- 2250
        b"010011000110_111100000000_000000100001_111110000000_000000000000_111000000000",	-- 2251
        b"010001101100_010101000000_000000100001_110011100110_010010110100_111000000000",	-- 2252
        b"010010000101_110100010000_000000100001_101110000000_000000000000_111011100000",	-- 2253
        b"010001101100_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 2254
        b"010001101101_110000010000_000000100001_111110000000_000000000000_111000000000",	-- 2255
        b"110000100000_010100000000_000001101001_110011000010_010010111001_111000000000",	-- 2256
        b"010010000101_110100010000_000000100001_100001000001_100110110010_111011100000",	-- 2257
        b"010001101101_110100010000_000000100001_110001000001_100111001001_111000000000",	-- 2260
        b"110000100100_010101000000_101110100001_011110000000_000000000000_111000000000",	-- 2261
        b"010000110101_111101100010_000001011101_110011000011_100001010111_111000000000",	-- 2262
        b"110001101101_110000000000_000000100001_110011000001_010010101111_111010000000",	-- 2263
        b"010010000101_110100010000_000000100001_100001000001_010100001111_111011100000",	-- 2264
        b"010001101101_110100010000_000000100001_110001000001_010100001011_111000000000",	-- 2265
        b"110000100100_010101000000_101110100001_011110000000_000000000000_111000000000",	-- 2266
        b"010000110101_111101100010_000001011101_110011000011_100001010111_111000000000",	-- 2267
        b"110001101101_110000000000_000000100001_110011000001_010010101111_111010000000",	-- 2270
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2271
        b"010001101101_110100010000_000000100001_110001000001_100111001001_111000000000",	-- 2272
        b"110010000000_000000000000_000000100001_100011000001_010010111110_111000000000",	-- 2273
        b"010000110101_111101100010_000000100001_110001010001_100001101100_111010000000",	-- 2274
        b"011101101100_010100000011_111110100001_110001000001_100111001010_111000000000",	-- 2275
        b"110000100101_010100000000_101111111101_110110000011_101000000000_111000000000",	-- 2276
        b"110010000000_000000000000_011000100001_100011000001_001100010000_111000000000",	-- 2277
        b"010001101101_110101110010_000000100001_111110000000_000000000000_111000000000",	-- 2300
        b"010000110101_111101100000_000000100001_010110000001_101000000000_111000000000",	-- 2301
        b"100101101011_010000000000_010010100001_110011000110_010110100111_111000000000",	-- 2302
        b"100100110000_010000000000_010010100001_110001000001_011000110111_111000000000",	-- 2303
        b"010011000110_111011100001_111110100001_110110000001_111100000000_111000000000",	-- 2304
        b"010001101011_010100100000_000000100001_110001000001_001100100111_111000000000",	-- 2305
        b"110010000000_000000000000_000000100001_100011010110_001110011111_111000000000",	-- 2306
        b"010001101100_010011110000_000000100001_111110000000_000000000000_111000000000",	-- 2307
        b"000101101100_111000000000_000010100001_110011011111_010011001101_111000000000",	-- 2310
        b"010011110000_010100100000_000000100001_111110000000_000000000000_111000000000",	-- 2311
        b"000101101000_010000100000_000010100001_111110000000_000000000000_111000000000",	-- 2312
        b"010010010000_011000100000_000000100001_111110000000_000000000000_111000000000",	-- 2313
        b"010010010000_110100100000_000000100001_111110000000_000000000000_111000000000",	-- 2314
        b"011000110100_110100100000_000110100001_101110000000_000000010111_111000100000",	-- 2315
        b"110011001100_111000000000_100000100001_010001100101_010011011010_111000000000",	-- 2316
        b"011101101100_110000100000_000001001001_100001000011_010011010010_111010000000",	-- 2317
        b"010010011000_110000011000_000000100001_111110000000_000000000000_111000000000",	-- 2320
        b"110010000000_000000000000_011000100001_101011000001_100001011000_111000000000",	-- 2321
        b"110010000000_000000000000_101000100001_101010000001_000000000000_111000000000",	-- 2322
        b"110010000000_000000000000_000000100001_100001011110_011000111010_111000000000",	-- 2323
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 2324
        b"010001101100_010011100000_000000100001_111011000001_001001110110_111000000000",	-- 2325
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2326
        b"010001101100_110101100000_000000100001_110001000001_100110110000_111000000000",	-- 2327
        b"010001101100_110011100000_000000100001_110001100101_010011011010_111000000000",	-- 2330
        b"010001101101_110100100000_000000100001_111011000001_010011001000_111000000000",	-- 2331
        b"110010000000_000000000000_000000100001_101010100001_000000000000_111000000000",	-- 2332
        b"010010001000_000011101000_000000100001_111010000001_000000000000_111000000000",	-- 2333
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2334
        b"010001101100_110101100000_000000100001_110001000001_100110110000_111000000000",	-- 2335
        b"110010000000_000000000000_000000100001_100001000001_010011101100_111000000000",	-- 2336
        b"010001101100_110011100000_000000100001_110001100101_010011011010_111000000000",	-- 2337
        b"010001101101_110100100000_000000100001_110011000001_010011001101_111000000000",	-- 2340
        b"110010000000_000000000000_000000100001_100001011110_011000111010_111000000000",	-- 2341
        b"010001101000_011100100000_000000100001_110001000001_100111001001_111000000000",	-- 2342
        b"010001101011_110100100000_000000100001_110001000001_100111001000_111000000000",	-- 2343
        b"110010000000_000000000000_000000100001_100001000001_100110110000_111000000000",	-- 2344
        b"010001101100_110101100000_000000100001_110001000001_100110110000_111000000000",	-- 2345
        b"010001101100_110011100000_000000100001_110001100101_010011011010_111000000000",	-- 2346
        b"010001101101_110100100000_000000100001_110011000001_010011001101_111000000000",	-- 2347
        b"110010000000_000000000000_000000100001_100001000001_010011101100_111000000000",	-- 2350
        b"010001101100_010011100000_011000100001_111011000001_001100010000_111000000000",	-- 2351
        b"010001101100_110101100000_000000100001_110011010110_001110011111_111000000000",	-- 2352
        b"010001101100_010100100000_000000100001_111011000001_010011011110_111000000000",	-- 2353
        b"110010000000_000000000000_000110100001_101110000000_000101101111_111000100000",	-- 2354
        b"010010001000_000000100000_000000100001_101110000000_000001000000_111000100000",	-- 2355
        b"011101101000_110000100000_000000100001_000001011110_011000111010_111010000000",	-- 2356
        b"110010000000_000000000000_000001001001_101010000010_000000000000_111000000000",	-- 2357
        b"010111001000_110000000001_010011101001_110011000010_010011110000_111000000000",	-- 2360
        b"100111001111_111000000001_010010100001_111110000000_000000000000_111000000000",	-- 2361
        b"010010010000_010000100000_000001101001_110011000011_010011110100_111010000000",	-- 2362
        b"010010001000_000100011001_001100100001_111010000001_000000000000_111000000000",	-- 2363
        b"010111001000_110000000001_010010100001_011110000000_000000000000_111000000000",	-- 2364
        b"010000110111_111100011001_001101001001_110011000010_010011110100_111000000000",	-- 2365
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 2366
        b"110010000000_000000000000_000000100001_100011010110_010011111001_111000000000",	-- 2367
        b"110010000000_000000000000_000000100001_100001011110_011000111010_111000000000",	-- 2370
        b"010001101000_011101100000_000000100001_110011000001_100011111001_111000000000",	-- 2371
        b"010010001000_000000000000_000001001001_110011000010_010011111110_111000000000",	-- 2372
        b"010001101100_010011100000_000001011101_110011000010_010011111110_111000000000",	-- 2373
        b"010000110101_110101100000_000000100001_011110000000_000000000000_111000000000",	-- 2374
        b"010001101000_010000000010_000001011101_110011000011_010011111100_111000000000",	-- 2375
        b"110010000000_000000000000_101110100001_101110000000_000000010000_111000000000",	-- 2376
        b"110011000111_111000000000_000000100001_111011000001_001100010000_111010000000",	-- 2377
        b"110010000000_000000000000_000110100001_101110000000_000000100000_111000100000",	-- 2400
        b"100101101011_010000000000_010010100001_111100000000_000000000011_111000000000",	-- 2401
        b"100100110000_010000000000_010010100001_111001000000_010100000010_111000000000",	-- 2402
        b"010010000000_000000100000_000000100001_100001000001_011001011100_111010000000",	-- 2403
        b"110011000000_010000011000_011001101001_111011000010_001100010000_111000000000",	-- 2404
        b"010010010000_010000011000_000000100001_110011000001_010110100111_111000000000",	-- 2405
        b"011011000111_110011000000_000000100001_100011011110_001100011101_111000000000",	-- 2406
        b"010011001111_111110000000_000000100001_110011000110_001100011101_111000000000",	-- 2407
        b"010001101101_110011000001_101000100001_111011000001_001100100001_111100100000",	-- 2410
        b"010010001000_000110010000_000000100001_101110000000_000000100000_111000100000",	-- 2411
        b"110010000000_000000000000_000000100001_100011000001_010100001100_111000000000",	-- 2412
        b"010010001000_000110010000_000000100001_101110000000_000010000000_111000100000",	-- 2413
        b"110010000000_000000000000_000000100001_100001000001_010100011010_111000000000",	-- 2414
        b"011111000110_111100000001_111110100001_110001000001_100111001001_111000000000",	-- 2415
        b"110010000000_000000000000_000000100001_100011000001_010100010100_111000000000",	-- 2416
        b"010010001000_000110010000_000000100001_101110000000_000000100000_111000100000",	-- 2417
        b"110010000000_000000000000_000000100001_100011000001_010100010010_111000000000",	-- 2420
        b"010010001000_000110010000_000000100001_101110000000_000010000000_111000100000",	-- 2421
        b"110010000000_000000000000_000000100001_100001000001_010100011010_111000000000",	-- 2422
        b"011111000110_111100000001_111110100001_110001000001_100110110011_111000000000",	-- 2423
        b"110010000000_000000000000_000110100001_101110000000_000101110010_111000100000",	-- 2424
        b"010010000000_000000101000_100000100001_101110000000_000000000000_111010000000",	-- 2425
        b"110010000000_000000000000_000110100001_101110000000_000101110011_111000100000",	-- 2426
        b"010010000000_000000110000_000000100001_101110000000_000000000000_111010000000",	-- 2427
        b"110001101000_110000000000_000000100001_111110000000_000000000000_111100000000",	-- 2430
        b"110011000111_111000100000_000000100001_111010000001_000000000000_111010000000",	-- 2431
        b"010010000110_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 2432
        b"110011000000_010110000000_000001101001_111010000010_000000000000_111000000000",	-- 2433
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 2434
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 2435
        b"110011000000_010000011000_000000100001_011110000000_000000000000_111000000000",	-- 2436
        b"110010000000_000000000000_000110100001_101110000000_000101110011_111000100000",	-- 2437
        b"010010000000_000000000000_000001001001_100001000011_010011010010_111010000000",	-- 2440
        b"100100110000_010000001000_010010100001_111110000000_000000000000_111000000000",	-- 2441
        b"100101101000_010000001000_010010100001_111110000000_000000000000_111000000000",	-- 2442
        b"110011000111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 2443
        b"110001101000_010000000000_000000100001_111010000001_000000000000_111100000000",	-- 2444
        b"010011000110_111100000001_111110100001_110001011110_011000111010_111000000000",	-- 2445
        b"010010001000_000000000000_000000100001_101110000000_010100101001_111000100000",	-- 2446
        b"110010000000_000000000000_000000100001_100001000001_101000001111_111000000000",	-- 2447
        b"010010001000_000000000000_000000010100_110001100000_100100010110_111000000000",	-- 2450
        b"010011000111_010100000000_101110100001_111110000000_000000000000_111000000000",	-- 2451
        b"010010001000_000000100000_000000100001_101110000000_001000000000_111000100000",	-- 2452
        b"010010000000_110000100000_000000100001_100001100000_011001100000_111011100000",	-- 2453
        b"010011110100_010000000000_011000100001_111011000001_001100010000_111010000000",	-- 2454
        b"110011000111_011101000000_101110100001_010110010111_101100000000_111000000000",	-- 2455
        b"110010000000_000000000000_011001000001_100011000010_010100110001_111000000000",	-- 2456
        b"010000110101_010101100000_000000100001_110011101111_100011100011_111010000000",	-- 2457
        b"010000110111_110101100000_000000100001_110011000001_100011100011_111010000000",	-- 2460
        b"010000110101_110101010000_011000100001_111110000000_000000000000_111000000000",	-- 2461
        b"010010000101_110101100000_000000100001_101110000000_000000000000_111011100000",	-- 2462
        b"010000110101_110101000000_000000011101_110011000011_001100010000_111010000000",	-- 2463
        b"110001101101_110000000000_000000011101_110001000010_100001100111_111000000000",	-- 2464
        b"110010000000_000000000000_000000100001_100011000001_100001011000_111000000000",	-- 2465
        b"010001101100_010001011000_000000100001_111110000000_000000000000_111000000000",	-- 2466
        b"011001101000_011000000000_000110100001_101110000000_000001100101_111000100000",	-- 2467
        b"010010000000_000010100000_000000100001_100011010111_010101000000_111010000000",	-- 2470
        b"110011000111_011101100000_000000100001_011110000000_000000000000_111000000000",	-- 2471
        b"010010000111_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 2472
        b"010011000000_010100101000_000001000001_110011000010_010101000001_111000000000",	-- 2473
        b"010001101101_110101100010_010000100001_111110000000_000000000000_111000000000",	-- 2474
        b"011101101101_110100000001_111110100001_110001000001_100111001010_111000000000",	-- 2475
        b"010010010010_110000011000_101110100001_111110000000_000000000000_111000000000",	-- 2476
        b"010001101001_011011100000_000000100001_110011000001_100011100011_111000000000",	-- 2477
        b"010011001111_111100101000_000000100001_111110000000_000000000000_111000000000",	-- 2500
        b"010000110101_111101101000_000000100001_111110000000_000000000000_111000000000",	-- 2501
        b"010001101101_110101110010_000000100001_111110000000_000000000000_111000000000",	-- 2502
        b"010001101101_110100010000_011000100001_110001000001_100111001001_111000000000",	-- 2503
        b"110011000111_110101100000_101110100001_011110000000_000000000000_111000000000",	-- 2504
        b"010010010010_110000011000_000000100001_111110000000_000000000000_111000000000",	-- 2505
        b"010001101001_011011100000_011001001001_111011000011_100011100011_111000000000",	-- 2506
        b"110001101101_110000000000_000000100001_110011000001_010101010110_111010000000",	-- 2507
        b"010001101011_110100100001_111110100001_110110000001_101000000000_111000000000",	-- 2510
        b"110001101011_110000000001_111110100001_111110000000_000000000000_111000000000",	-- 2511
        b"110011000111_011101000000_000000100001_010011010111_010101010000_111000000000",	-- 2512
        b"110010000000_000000000000_000001000001_100011000010_010101010000_111000000000",	-- 2513
        b"010001101101_010100000010_000000100001_110001100110_010100001001_111000000000",	-- 2514
        b"011111000110_111100000001_111110100001_110001100111_100111001010_111000000000",	-- 2515
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 2516
        b"110001101101_010000000010_010000100001_111011000001_001100010000_111010000000",	-- 2517
        b"010000110101_111101001000_000000100001_111110000000_000000000000_111000000000",	-- 2520
        b"010001101101_010101010010_000000100001_111110000000_000000000000_111000000000",	-- 2521
        b"010001101101_010100010000_000000100001_110001100110_010100001001_111000000000",	-- 2522
        b"011111000110_111100000001_111110100001_110001100111_100111001010_111000000000",	-- 2523
        b"110011000111_110101000000_101110100001_011110000000_000000000000_111000000000",	-- 2524
        b"110011000111_111101000000_011001001001_111011000011_001100010000_111010000000",	-- 2525
        b"110010000000_000000000000_000000100001_100001000001_100001100111_111000000000",	-- 2526
        b"110010000000_000000000000_011000100001_101011000001_100001011000_111000000000",	-- 2527
        b"110011000111_011101100000_000000100001_010011010111_010101100111_111000000000",	-- 2530
        b"010001101100_010010100000_000001000001_110011000010_010101101000_111000000000",	-- 2531
        b"011101101101_110100000000_000000100001_110011011101_010101011110_111000000000",	-- 2532
        b"010011000110_111100000000_010000100001_110001100110_010100001111_111000000000",	-- 2533
        b"011101101100_010100000001_111110100001_110001100111_100110110011_111000000000",	-- 2534
        b"110010000000_000000000000_011000100001_100011000001_010101100000_111000000000",	-- 2535
        b"010011000110_111100000000_000000100001_110001100110_010100001111_111000000000",	-- 2536
        b"011101101100_010100000001_111110100001_110001100111_100110110011_111000000000",	-- 2537
        b"010001101010_110100000000_000000100001_110001100110_010100001011_111000000000",	-- 2540
        b"011111000110_111100000001_111110100001_110001100111_100111001010_111000000000",	-- 2541
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 2542
        b"110000110111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2543
        b"010001101101_110100010000_011000100001_110001100110_010100001111_111000000000",	-- 2544
        b"011111000110_111100000001_111110100001_110001100111_100110110011_111000000000",	-- 2545
        b"110010000000_000000000000_010000100001_100011000001_010101101011_111000000000",	-- 2546
        b"010001101100_010010100000_000000100001_111110000000_000000000000_111000000000",	-- 2547
        b"010001101011_110100000000_000000100001_110011011101_010101100100_111000000000",	-- 2550
        b"010001101101_110100010000_011000100001_110001100110_010100001111_111000000000",	-- 2551
        b"011111000110_111100000001_111110100001_110001100111_100110110011_111000000000",	-- 2552
        b"010001101010_110100000000_000000100001_110001100110_010100001011_111000000000",	-- 2553
        b"011111000110_111100000001_111110100001_110001100111_100111001010_111000000000",	-- 2554
        b"110011000111_110101100000_000000100001_011110000000_000000000000_111000000000",	-- 2555
        b"010000010101_111101100010_101110100001_111110000000_000000000000_111000000000",	-- 2556
        b"010000110111_111101110000_011001001001_111011000011_100011100011_111000000000",	-- 2557
        b"110011000111_111101100000_000000100001_110011000001_010101010110_111010000000",	-- 2560
        b"110010010111_110011000000_000001101001_110011000011_001110011111_111000000000",	-- 2561
        b"110011000111_011101100000_000000100001_010011010110_010101110101_111000000000",	-- 2562
        b"010001101101_110100010000_000000100001_110001000001_100110110010_111000000000",	-- 2563
        b"010001101100_110011110000_000000100001_110011000001_010101101101_111000000000",	-- 2564
        b"010001101101_110100010000_011001000001_110011000011_010101111000_111000000000",	-- 2565
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2566
        b"010001101100_110011100000_000000100001_110011000001_010101101101_111000000000",	-- 2567
        b"010001101101_110100000000_010000100001_110001000001_100110110010_111000000000",	-- 2570
        b"010001101100_110011100000_101110100001_111110000000_000000000000_111000000000",	-- 2571
        b"110000110111_111101100000_011000100001_111011000001_001100010000_111010000000",	-- 2572
        b"110010000000_000000000000_000110100001_101110000000_000001100101_111000100000",	-- 2573
        b"010010000000_000010000000_000000100001_100011010111_010101111110_111010000000",	-- 2574
        b"010011000110_111100100000_101110100001_110110000001_100100000000_111000000000",	-- 2575
        b"010001101000_011100101000_101110100001_110110000001_100100000000_111000000000",	-- 2576
        b"110010000000_000000000000_000000100001_100011000111_001110011111_111000000000",	-- 2577
        b"110010000000_000000000000_000000100001_100001000001_100111001001_111000000000",	-- 2600
        b"010001101100_010100010010_000000100001_111110000000_000000000000_111000000000",	-- 2601
        b"010010010010_010000011000_000000100001_111110000000_000000000000_111000000000",	-- 2602
        b"010001101100_010011100000_011000100001_111011000001_001100010000_111000000000",	-- 2603
        b"110011000111_111100100000_000000100001_110011000001_010110000010_111010000000",	-- 2604
        b"010001101101_110100100000_000000100001_110001000001_100111001001_111000000000",	-- 2605
        b"010010000100_010101100000_000000100001_101110000000_000000000000_111011100000",	-- 2606
        b"010001101011_110101110000_000000100001_111110000000_000000000000_111000000000",	-- 2607
        b"010001101100_010011100000_000000100001_111110000000_000000000000_111000000000",	-- 2610
        b"010001101011_110011110010_000000100001_110011000001_100011100010_111000000000",	-- 2611
        b"010001101100_010010100000_000000100001_111110000000_000000000000_111000000000",	-- 2612
        b"010010000101_110100010000_000000100001_100001000001_100110110010_111011100000",	-- 2613
        b"010001101010_110011100000_101110100001_111110000000_000000000000_111000000000",	-- 2614
        b"110001101100_110000000000_011000100001_110011000001_001100010000_111010000000",	-- 2615
        b"110000100101_010101100000_000000100001_010110000001_101000000000_111000000000",	-- 2616
        b"010001101101_110101100010_000001101000_110011000010_010000111101_111000000000",	-- 2617
        b"110010000000_000000000000_000001001101_100110000011_101000000000_111000000000",	-- 2620
        b"110010000000_000000000000_000000100001_100011000001_010000111000_111000000000",	-- 2621
        b"010000110111_111101100000_000001001001_010110000010_101000000000_111000000000",	-- 2622
        b"110010000000_000000000000_000001001101_100011000011_010000111101_111000000000",	-- 2623
        b"110010000000_000000000000_000000100001_100011000001_010001000000_111000000000",	-- 2624
        b"110010000000_000000000000_000001000101_100110000011_101100000000_111000000000",	-- 2625
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2626
        b"110010000000_000000000000_000001001001_100110000011_101100000000_111000000000",	-- 2627
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2630
        b"110010000000_000000000000_000001000001_100110000011_101100000000_111000000000",	-- 2631
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2632
        b"110010000000_000000000000_000001000101_100110000010_101100000000_111000000000",	-- 2633
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2634
        b"110010000000_000000000000_000001001001_100110000010_101100000000_111000000000",	-- 2635
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2636
        b"110010000000_000000000000_000001000001_100110000010_101100000000_111000000000",	-- 2637
        b"010001101011_110011110010_000000100001_110110000001_101100000000_111000000000",	-- 2640
        b"110010000000_000000000000_011001011101_100110000011_101100000000_111000000000",	-- 2641
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2642
        b"110010000000_000000000000_011001001001_100110000011_101100000000_111000000000",	-- 2643
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2644
        b"110010000000_000000000000_011001000001_100110000011_101100000000_111000000000",	-- 2645
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2646
        b"010001101100_010011100000_011000100001_110110000001_101100000000_111000000000",	-- 2647
        b"110010000000_000000000000_011001011111_100110000011_101100000000_111000000000",	-- 2650
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2651
        b"110010000000_000000000000_011001001001_100110000010_101100000000_111000000000",	-- 2652
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2653
        b"110010000000_000000000000_011001000001_100110000010_101100000000_111000000000",	-- 2654
        b"010001101100_010011100000_000000100001_110110000001_101100000000_111000000000",	-- 2655
        b"110010000000_000000000000_011000100001_101011000110_001100010000_111000000000",	-- 2656
        b"110011000111_111101100000_000000100001_111011000001_001100010000_111010000000",	-- 2657
        b"010010001000_000101100000_000000100001_110110000001_100100000000_111000000000",	-- 2660
        b"010011000101_010101100000_000000100001_110110000001_101000000000_111000000000",	-- 2661
        b"010010010101_010101100000_000000100001_110110000001_101000000000_111000000000",	-- 2662
        b"110010000000_000000000000_000000100001_100001000001_001110011000_111000000000",	-- 2663
        b"110010000000_000000000000_101110100001_100110000001_101000000000_111000000000",	-- 2664
        b"010001110101_110101100000_000000100001_110011000001_010110110001_111000000000",	-- 2665
        b"010010110101_010101100000_000000100001_111110000000_000000000000_111000000000",	-- 2666
        b"110010000000_000000000000_000000100001_100110000001_101000000000_111000000000",	-- 2667
        b"010011110101_010101100000_000000100001_110110000001_101000000000_111000000000",	-- 2670
        b"010001110101_110101100000_000000100001_111110000000_000000000000_111000000000",	-- 2671
        b"010010010101_010101100000_000000100001_110110000001_101000000000_111000000000",	-- 2672
        b"010010100101_010101100000_000000100001_110110000001_101000000000_111000000000",	-- 2673
        b"010001110101_110101100000_000000100001_110110000001_101000000000_111000000000",	-- 2674
        b"010001110101_010101000000_000000100001_110011000001_010110111000_111000000000",	-- 2675
        b"010001110101_110101100000_000000100001_110110000001_101000000000_111000000000",	-- 2676
        b"010001110101_110101100000_000000100001_110011000001_010110111000_111000000000",	-- 2677
        b"110011000101_010101100000_000000100001_100011000001_010110111110_111000000000",	-- 2700
        b"010000001000_000101100000_000000100001_110110000001_100100000000_111000000000",	-- 2701
        b"010001101101_010101110000_000000100001_110110000001_101000000000_111000000000",	-- 2702
        b"010001101100_010101101001_111110100001_111110000000_000000000000_111000000000",	-- 2703
        b"010011000110_111101100000_000000100001_110011010010_100011100010_111000000000",	-- 2704
        b"110001101011_110000000001_111110100001_110011011101_100011100010_111000000000",	-- 2705
        b"110010000000_000000000000_101110100001_100110010111_101000000000_111000000000",	-- 2706
        b"010001101101_111101101000_000000100001_110011000001_100011100011_111000000000",	-- 2707
        b"010010000101_010101000000_000000100001_101110000000_000000000000_111011100000",	-- 2710
        b"010001101101_010101101000_000000100001_110110000001_101000000000_111000000000",	-- 2711
        b"010010000101_110101001000_000000100001_100110000001_101000000000_111011100000",	-- 2712
        b"010010000101_110101101000_000000100001_100110000001_101000000000_111011100000",	-- 2713
        b"010011000111_110101100000_000000100001_110110000001_101100000000_111000000000",	-- 2714
        b"110001101101_110000000000_000000100001_011110000000_000000000000_111000000000",	-- 2715
        b"010010001000_000101110000_000001011101_110110000011_101100000000_111000000000",	-- 2716
        b"010000001000_000101110000_000000100001_110110000001_101100000000_111000000000",	-- 2717
        b"010001101101_010101101000_000000100001_110110000001_101000000000_111000000000",	-- 2720
        b"010010000101_010101000000_000000100001_101110000000_000000000000_111011100000",	-- 2721
        b"010001101101_010101110000_000000100001_110110000001_101000000000_111000000000",	-- 2722
        b"010010000101_110101010000_000000100001_100110000001_101000000000_111011100000",	-- 2723
        b"010010000101_110101110000_000000100001_100011000001_100011101101_111011100000",	-- 2724
        b"010010001000_000101101000_000000100001_110110000001_101100000000_111000000000",	-- 2725
        b"010010010111_110101100000_000000100001_110110101111_101100000000_111000000000",	-- 2726
        b"010000001000_000101101000_000000100001_110110000001_101100000000_111000000000",	-- 2727
        b"010010001000_000100001000_000000100001_110011000001_010111011101_111000000000",	-- 2730
        b"010010001000_000100001000_000000100001_111110000000_000000000000_111000000000",	-- 2731
        b"010010000100_010100000000_000000100001_100011000001_010111011101_111011100000",	-- 2732
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2733
        b"010001101100_110100000000_101110100001_111110000000_000000000000_111000000000",	-- 2734
        b"010010000000_000101100000_011000100001_100110000001_100100000000_111010000000",	-- 2735
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2736
        b"010010000100_110100000000_101110100001_101110000000_000000000000_111011100000",	-- 2737
        b"010010000000_000101100000_011000100001_100110000001_100100000000_111010000000",	-- 2740
        b"110011000100_010101100000_000001101001_110110000011_101000000000_111000000000",	-- 2741
        b"010001101011_110011110010_000000100001_110110000001_101000000000_111000000000",	-- 2742
        b"110011000100_010101100000_000001101001_110110000010_101000000000_111000000000",	-- 2743
        b"010001101011_110011110010_000000100001_110110000001_101000000000_111000000000",	-- 2744
        b"110010010100_010101100000_000000100001_111011000001_001100010000_111010000000",	-- 2745
        b"110010110100_010101100000_000000100001_111011000001_001100010000_111010000000",	-- 2746
        b"110011110100_010101100000_000000100001_111011000001_001100010000_111010000000",	-- 2747
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2750
        b"110010000000_000000000000_000000100001_100001000001_001100100111_111000000000",	-- 2751
        b"010010001000_000000000000_000000100001_101110000000_000100000000_111000100000",	-- 2752
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 2753
        b"011001101000_010000000000_000000100001_101110000000_000000000000_111000000000",	-- 2754
        b"010111001011_010000000000_000010100001_011110000000_000000000000_111000000000",	-- 2755
        b"010111001011_010000000000_000011001001_010011000010_010111111100_111000000000",	-- 2756
        b"010111001011_010000000000_000011001001_010011000011_010111110101_111000000000",	-- 2757
        b"010001101100_010000100000_000000100001_111110000000_000000000000_111000000000",	-- 2760
        b"100101101000_110000100000_010011101001_110001000011_010111110100_111000000000",	-- 2761
        b"100101101000_110000100000_010011101001_110001000011_010111110100_111000000000",	-- 2762
        b"110011000000_011100111000_000000100001_101110000000_000000000000_111000000000",	-- 2763
        b"010001101000_110000100010_000000100001_111010000001_000000000000_111000000000",	-- 2764
        b"010111001011_010000000000_000011001001_010011000011_001110011111_111000000000",	-- 2765
        b"010001101100_010001000000_000001001001_110011000011_010111111100_111000000000",	-- 2766
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 2767
        b"110010000000_000000000000_000110100001_101110000000_000000100000_111000100000",	-- 2770
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 2771
        b"110010010000_010100100000_000000100001_011110000000_000000000000_111000000000",	-- 2772
        b"010001101100_110000100000_000001001001_110011000011_001110011111_111000000000",	-- 2773
        b"110010000000_000000000000_000000100001_100110000001_100100000000_111000000000",	-- 2774
        b"110011000100_111000011000_000000100001_101110000000_000000000000_111000000000",	-- 2775
        b"000110001000_000010100000_001010100001_101110000000_000000000000_111000100000",	-- 2776
        b"000101101010_110010100000_000010100001_111110000000_000000000000_111000000000",	-- 2777
        b"000101101010_110010100000_000010100001_111110000000_000000000000_111000000000",	-- 3000
        b"110010000000_000000000000_000000100001_100001000001_011000001111_111000000000",	-- 3001
        b"110010000000_000000000000_000000100001_100001000001_011000011101_111000000000",	-- 3002
        b"010000110111_111010100000_000001101001_110011000011_011000000001_111000000000",	-- 3003
        b"110010000000_000000000000_000000100001_101011000001_001100010000_111000000000",	-- 3004
        b"110010000000_000000000000_000000100001_100001000001_011000001111_111000000000",	-- 3005
        b"110010000000_000000000000_000110100001_101110000000_000100100110_111000100000",	-- 3006
        b"110011000111_010000000000_000000100001_110001000001_011000011101_111010000000",	-- 3007
        b"011011000111_010000000000_000110100001_101110000000_000100100110_111000100000",	-- 3010
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3011
        b"110000011000_010000000010_000001101000_110011000011_011000001101_111000000000",	-- 3012
        b"010000110111_111010100000_000001101001_110011000011_011000000101_111000000000",	-- 3013
        b"110010000000_000000000000_000000100001_101011000001_001100010000_111000000000",	-- 3014
        b"110010000000_000000000000_000001011101_100011000010_011000001110_111000000000",	-- 3015
        b"110010000000_000000000000_000000100001_101011000001_001100010000_111000000000",	-- 3016
        b"010001101000_110000100010_000001111101_010011000010_011000011100_111000000000",	-- 3017
        b"000101101000_110100000000_010010100001_111110000000_000000000000_111000000000",	-- 3020
        b"000101101000_110100000000_010011010101_110011000010_011000011010_111000000000",	-- 3021
        b"110010000000_000000000000_000001010101_100011000010_011000010111_111000000000",	-- 3022
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3023
        b"010001101100_110001000000_000000100001_111100000000_000000000010_111000000000",	-- 3024
        b"010010000001_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3025
        b"100101101000_010000000000_010010100001_110011000001_011000011000_111000000000",	-- 3026
        b"100101101001_010000000000_010010100001_111100000000_000000000011_111000000000",	-- 3027
        b"100100110000_010000000000_010010100001_111001000000_011000011000_111000000000",	-- 3030
        b"010010000000_010000000000_000000100001_101010000001_000000000000_111011100000",	-- 3031
        b"010001101001_010000000000_000001010101_111010000010_000000000000_111000000000",	-- 3032
        b"010010000000_010000000000_000000100001_101010000001_000000000000_111011100000",	-- 3033
        b"010001101001_010000000000_000000100001_111010000001_000000000000_111000000000",	-- 3034
        b"010001101001_110001100010_000000100001_111110000000_000000000000_111000000000",	-- 3035
        b"000101101001_110100000000_010010100001_111110000000_000000000000_111000000000",	-- 3036
        b"000101101001_110100000000_010011010101_110011000010_011000101010_111000000000",	-- 3037
        b"110010000000_000000000000_000001010101_100011000010_011000100110_111000000000",	-- 3040
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3041
        b"010001101100_110010000000_000000100001_111100000000_000000000011_111000000000",	-- 3042
        b"110010000000_000000000000_000110100001_101110000000_000100101100_111000100000",	-- 3043
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3044
        b"100101101000_010000000000_010010100001_110011000001_011000101000_111000000000",	-- 3045
        b"110010000000_000000000000_000110100001_101110000000_000100101101_111000100000",	-- 3046
        b"100101101010_010000000000_010010100001_111100000000_000000000011_111000000000",	-- 3047
        b"100100110000_010000000000_010010100001_111001000000_011000101000_111000000000",	-- 3050
        b"010010000000_000100100000_000000100001_101010000001_000000000000_111010000000",	-- 3051
        b"010010000111_010100100000_000001010101_100011000010_011000101111_111011100000",	-- 3052
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3053
        b"010010010100_110010000000_000000100001_111110000000_000000000000_111000000000",	-- 3054
        b"010011000100_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 3055
        b"010011110000_010010000000_000000100001_111010000001_000000000000_111000000000",	-- 3056
        b"011010010111_010010000000_000000100001_101110000000_000000000000_111000000000",	-- 3057
        b"010011000111_010000000000_000000100001_111110000000_000000000000_111000000000",	-- 3060
        b"010011111000_010100100000_000000100001_110001000001_100111001001_111000000000",	-- 3061
        b"011101101100_010100000011_111110100001_110001000001_100110110011_111000000000",	-- 3062
        b"010001101100_110010000000_000000100001_111010000001_000000000000_111000000000",	-- 3063
        b"100101101011_010000000000_010010100001_110001011110_011000111010_111000000000",	-- 3064
        b"100100110000_010000000000_010010100001_110001000001_011000110111_111000000000",	-- 3065
        b"110010000000_000000000000_000000100001_100110000001_111000000000_111000000000",	-- 3066
        b"100101101000_010000000000_010010100001_111010000001_000000000000_111100100000",	-- 3067
        b"110010000000_000000000000_000000100001_100001011110_011000111010_111000000000",	-- 3070
        b"110010000000_000000000000_000000100001_101011000001_001100010000_111000000000",	-- 3071
        b"010010001000_000000000000_000000100001_101010011111_100000000000_111000100000",	-- 3072
        b"010010000000_010000000000_000000100001_101010100110_000000000000_111011100000",	-- 3073
        b"110011000000_010000011000_000001101001_111010000011_000000000000_111000000000",	-- 3074
        b"110010000000_000000000000_000000100001_101011000001_001110011111_111000000000",	-- 3075
        b"000101101101_111101100001_010010100001_101110000000_100000000010_111000100000",	-- 3076
        b"010010000101_110101100000_000000100001_100011000001_100011111001_111011100000",	-- 3077
        b"000101101101_111000000001_010010100001_101110000000_000000001000_111000100000",	-- 3100
        b"110011000000_010100000000_000001101001_110011000011_001110011111_111000000000",	-- 3101
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 3102
        b"011000110000_010000000000_000110100001_101110000000_000101101110_111000100000",	-- 3103
        b"010010001000_000000100000_000000100001_101110000000_111111110000_111000100000",	-- 3104
        b"010011000100_010000100000_000000100001_111110000000_000000000000_111000000000",	-- 3105
        b"010010000000_000000000000_000000100001_100001000001_011001011010_111010000000",	-- 3106
        b"010010000000_110000100000_000000100001_100001000001_011001011101_111011100000",	-- 3107
        b"010010001000_000000100000_000000100001_101110000000_000000000111_111000100000",	-- 3110
        b"010010010000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 3111
        b"010011000100_010000100000_000000100001_111110000000_000000000000_111000000000",	-- 3112
        b"110011110000_110000000000_000000100001_111110000000_000000000000_111010000000",	-- 3113
        b"110111001100_010000000000_010011101001_110001000011_011001001111_111000000000",	-- 3114
        b"110010000000_000000000000_000000100001_100001000001_011010010101_111000000000",	-- 3115
        b"110010000000_000000000000_011000100001_101011000001_001100010000_111000000000",	-- 3116
        b"110010000000_000000000000_000110100001_101110000000_000101101110_111000100000",	-- 3117
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 3120
        b"010010001000_000010100000_000110100001_101110000000_000010000000_111000100000",	-- 3121
        b"010010001000_000010100000_000000100001_101110000000_100010000000_111000100000",	-- 3122
        b"010010000010_010010000000_000000100001_101110000000_000000000000_111011100000",	-- 3123
        b"100100110010_010010000000_010010100001_111110000000_000000000000_111010000000",	-- 3124
        b"011001101010_110000000010_000000100001_101100000000_000000111101_111000000000",	-- 3125
        b"011001101000_000000000010_000110100001_111110000000_000000000000_111000000000",	-- 3126
        b"110010001000_000000000000_000000100001_111001000000_011001010110_111010000000",	-- 3127
        b"110010001000_000000000000_000000100001_110001000001_011010010101_111100000000",	-- 3130
        b"110010000000_000000000000_000000100001_100011000001_011101000000_111000000000",	-- 3131
        b"110111001100_010000000000_010011101001_110001000011_011001100000_111000000000",	-- 3132
        b"110111001100_010000000000_010011101001_111010000010_000000000000_111000000000",	-- 3133
        b"010010010000_110000000000_000000100001_111010000001_000000000000_111000000000",	-- 3134
        b"110111001100_010000000000_010011101001_110011000010_011001011111_111000000000",	-- 3135
        b"010010010000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 3136
        b"110111001100_010000000000_010011101001_111010000010_000000000000_111000000000",	-- 3137
        b"010011110000_110000000000_000000100001_111010000001_000000000000_111000000000",	-- 3140
        b"110010000000_000000000000_000000100001_100001000001_011001100011_111000000000",	-- 3141
        b"110010000000_000000000000_000000100001_100011000001_100011111001_111000000000",	-- 3142
        b"110010000000_000000000000_000110100001_101110000000_000101101110_111000100000",	-- 3143
        b"010010000000_000101100000_000000100001_101110000000_000000000000_111010000000",	-- 3144
        b"010010000101_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 3145
        b"110011000101_110000000000_000000100001_011110000000_000000000000_111000000000",	-- 3146
        b"010010001000_000000000000_000001001001_101010000010_000000001000_111000100000",	-- 3147
        b"010011110000_010101100000_000000100001_111010000001_000000000000_111000000000",	-- 3150
        b"110010000000_000000000000_000000100001_100001000001_011001100011_111000000000",	-- 3151
        b"010010001000_000101101000_000000100001_110011000001_011010111110_111000000000",	-- 3152
        b"110010000000_000000000000_000000100001_100001000001_011001100011_111000000000",	-- 3153
        b"010010001000_000101101000_000000100001_110011000001_011011000001_111000000000",	-- 3154
        b"010010001000_000000000000_000000100001_101110000000_111100000000_111000100000",	-- 3155
        b"100100110000_010000000000_010010100001_110001000001_011011010010_111000000000",	-- 3156
        b"000110001000_000000100000_001010100001_111110000000_000000000000_111000000000",	-- 3157
        b"010010001000_000001000000_000000100001_101110000000_000001111111_111000100000",	-- 3160
        b"011001101001_010000000010_000110100001_101110000000_000101110001_111000100000",	-- 3161
        b"010011000100_010001000000_000000100001_111110000000_000000000000_111000000000",	-- 3162
        b"010010000000_000000000000_000000100001_100001000001_011001011010_111010000000",	-- 3163
        b"010010001000_000000000000_000000100001_101110000000_111100000001_111000100000",	-- 3164
        b"100100110000_010000000000_010010100001_110001000001_011011010010_111000000000",	-- 3165
        b"000110001000_000000100000_001010100001_111110000000_000000000000_111000000000",	-- 3166
        b"010001101110_110001000000_000000100001_111110000000_000000000000_111000000000",	-- 3167
        b"011001101001_010000000010_000110100001_101110000000_000101110001_111000100000",	-- 3170
        b"010011000100_010001000000_000000100001_111110000000_000000000000_111000000000",	-- 3171
        b"101110000000_000000000000_110010100001_100001000001_011001011010_111010000000",	-- 3172
        b"010001101001_010000100000_000000100001_110001000001_011001011101_111000000000",	-- 3173
        b"110011000111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 3174
        b"110010000000_000000000000_000110100001_101110000000_000101110000_111000100000",	-- 3175
        b"110111001100_010000000000_010010100001_011110000000_000000000000_111000000000",	-- 3176
        b"010010000000_000000100000_000001001001_100011000010_011010000001_111010000000",	-- 3177
        b"010011110001_010000100000_000000100001_111110000000_000000000000_111010000000",	-- 3200
        b"110111001100_010000000000_010011101001_110011000010_011010000100_111000000000",	-- 3201
        b"110010000000_000000000000_000000100001_100001000001_011010001000_111000000000",	-- 3202
        b"110010000000_000000000000_011000100001_101011000001_001100010000_111000000000",	-- 3203
        b"110011001100_010000000000_000001101001_110011000010_011010000110_111000000000",	-- 3204
        b"010010010001_010000100000_000000100001_111110000000_000000000000_111010000000",	-- 3205
        b"110010000000_000000000000_000000100001_100001000001_011010010100_111000000000",	-- 3206
        b"110010000000_000000000000_011000100001_101011000001_001100010000_111000000000",	-- 3207
        b"110010000000_000000000000_000110100001_101110000000_000101101111_111000100000",	-- 3210
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 3211
        b"110010000000_000000000000_000110100001_101110000000_000101110000_111000100000",	-- 3212
        b"110010001000_000000000000_000100100001_111110000000_000000000000_111010000000",	-- 3213
        b"110010000000_000000000000_000110100001_101110000000_000101110001_111000100000",	-- 3214
        b"010010001000_000100011001_001100100001_110011000001_011010010100_111010000000",	-- 3215
        b"110010000000_000000000000_000110100001_101110000000_000101110001_111000100000",	-- 3216
        b"010010001000_000000100000_000000100001_101110000000_000011000000_111000100000",	-- 3217
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3220
        b"110001101000_010000000000_000001111101_110011000011_011010010011_111000000000",	-- 3221
        b"010011110000_010000100000_000000100001_111110000000_000000000000_111000000000",	-- 3222
        b"110001110000_110000000001_110100100001_111010000001_000000000000_111000000000",	-- 3223
        b"110010000000_000000000000_000000100001_100001000001_011010001110_111000000000",	-- 3224
        b"110010000000_000000000000_000110100001_101110000000_000101110000_111000100000",	-- 3225
        b"010010000000_000001100000_000000100001_101110000000_000000000000_111010000000",	-- 3226
        b"110010000000_000000000000_000110100001_101110000000_000101101110_111000100000",	-- 3227
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3230
        b"010010000000_010000100000_000000100001_101110000000_000000000000_111011100000",	-- 3231
        b"110011000000_010000100000_000001101001_110001000011_011010101001_111000000000",	-- 3232
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 3233
        b"100100110000_010000000000_010010100001_101110000000_010010010000_111000100000",	-- 3234
        b"011001101000_010000000000_000000100001_101100000000_000000000111_111000000000",	-- 3235
        b"010010001000_000001000000_000110100001_101110000000_000010000000_111000100000",	-- 3236
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3237
        b"100111001000_010000100000_010011101001_110011000010_011010100010_111000000000",	-- 3240
        b"110011000000_010000100000_000001101001_110001000011_011010101001_111000000000",	-- 3241
        b"010010001000_000000000000_000000100001_101110000000_000000001000_111000100000",	-- 3242
        b"010000110000_010001000000_000110100001_111001000000_011010011111_111000000000",	-- 3243
        b"110010000000_000000000000_000110100001_101110000000_000101110010_111000100000",	-- 3244
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 3245
        b"110010000000_000000000000_000110100001_101110000000_000101110011_111000100000",	-- 3246
        b"110011110001_110001000000_000000100001_111110000000_000000000000_111010000000",	-- 3247
        b"110011110001_110001000000_000000100001_111010000001_000000000000_111100000000",	-- 3250
        b"010010001000_000000100000_000000100001_101110000000_000000000111_111000100000",	-- 3251
        b"010011000000_110000000000_000001101001_111010000010_000000000000_111000000000",	-- 3252
        b"010010001000_000000100000_000000100001_101110000000_000001011100_111000100000",	-- 3253
        b"110000110000_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3254
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3255
        b"010011110000_010001100000_000000100001_111010000001_000000000000_111000000000",	-- 3256
        b"110010000000_000000000000_000000100001_100001000001_011010110011_111000000000",	-- 3257
        b"110010000000_000000000000_000110100001_101110000000_000101110000_111000100000",	-- 3260
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3261
        b"010010000000_010101101000_000000100001_100011000001_100011111001_111011100000",	-- 3262
        b"110010000000_000000000000_000110100001_101110000000_000101110001_111000100000",	-- 3263
        b"010010001000_000000000000_000000100001_101110000000_000001111111_111000100000",	-- 3264
        b"011101101000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 3265
        b"110010000000_000000000000_000110100001_101110000000_000101101111_111000100000",	-- 3266
        b"110001101000_010000000000_000000100001_011110000000_000000000000_111000000000",	-- 3267
        b"010011001000_010101100000_000001011101_110011000011_011010111010_111000000000",	-- 3270
        b"010000111101_110101100010_000000100001_111110000000_000000000000_111000000000",	-- 3271
        b"010010000000_000000000000_000000100001_100100000001_000000000011_111010000000",	-- 3272
        b"100100110000_010000000000_010010100001_111000000000_000000000000_111000000000",	-- 3273
        b"010011110000_010101100000_000000100001_111010000001_000000000000_111000000000",	-- 3274
        b"110010000000_000000000000_000000100001_100001000001_011010110011_111000000000",	-- 3275
        b"110011000101_110100000000_011001101001_111011000011_001100010000_111000000000",	-- 3276
        b"010001101011_110011110010_000000100001_111011000001_001100010000_111000000000",	-- 3277
        b"110010000000_000000000000_000000100001_100001000001_011010110011_111000000000",	-- 3300
        b"110011000101_110100000000_011001101001_111011000010_001100010000_111000000000",	-- 3301
        b"010001101011_110011110010_000000100001_111011000001_001100010000_111000000000",	-- 3302
        b"010010001000_000000000000_000000100001_101110000000_111000000000_111000100000",	-- 3303
        b"100100110000_010000000000_010010100001_110001000001_011011010010_111000000000",	-- 3304
        b"110010000000_000000000000_000000100001_100001000001_100100010000_111000000000",	-- 3305
        b"010001101100_010000000000_000000100001_110001000001_011011001110_111000000000",	-- 3306
        b"110010000000_000000000000_000110100001_101110000000_000001010110_111000100000",	-- 3307
        b"010011001000_110001111001_011000100001_111110000000_000000000000_111000000000",	-- 3310
        b"011101101100_010000100000_110000100001_101110000000_000000000000_111010000000",	-- 3311
        b"001111000000_110100000001_010011101001_110001000011_011011001101_111000000000",	-- 3312
        b"110011001000_110000000000_000001101001_110011000011_100001010111_111000000000",	-- 3313
        b"110010000000_000000000001_010000100001_100011000001_100001010111_111000000000",	-- 3314
        b"110010000000_000000000000_111000100001_101010000001_000000000000_111000000000",	-- 3315
        b"110010000000_000000000000_000110100001_101110000000_000000010110_111000100000",	-- 3316
        b"100101101000_010000000000_010010100001_110100000001_000000000011_111000000000",	-- 3317
        b"100100110000_010000000000_010010100001_111000000000_000000000000_111000000000",	-- 3320
        b"011101101000_010000100000_000000100001_101010000001_000000000000_111010000000",	-- 3321
        b"100100110000_010000000000_010010100001_111110000000_000000000000_111000000000",	-- 3322
        b"100100110000_010000000000_010010100001_111110000000_000000000000_111000000000",	-- 3323
        b"110011000000_010100000000_000001101001_111010000010_000000000000_111000000000",	-- 3324
        b"110010000000_000000000000_000000100001_100011000001_001110011111_111000000000",	-- 3325
        b"110010000000_000000000000_000110100001_101110000000_000001010110_111000100000",	-- 3326
        b"010001101001_111000000000_000000100001_110001000001_011011001111_111000000000",	-- 3327
        b"010010000000_010000000000_000000100001_100001100000_011001100000_111011100000",	-- 3330
        b"100101101000_110000100000_010010100001_110001100100_011001100000_111000000000",	-- 3331
        b"010001101000_010101100000_000000100001_110011000001_100011111001_111000000000",	-- 3332
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3333
        b"110010000000_000000000000_000000100001_100001000001_100100010000_111000000000",	-- 3334
        b"000110001000_000001000000_001010100001_111110000000_000000000000_111000000000",	-- 3335
        b"011001101001_010000000000_000110100001_101110000000_000101110010_111000100000",	-- 3336
        b"010111001100_110000000000_000010100001_011110000000_000000000000_111000000000",	-- 3337
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 3340
        b"010010001000_000000100000_000000100001_101110000000_111111000000_111000100000",	-- 3341
        b"010010000001_110001100000_000001001001_100011000010_011011100110_111011100000",	-- 3342
        b"010010010001_110001000000_000000100001_111110000000_000000000000_111000000000",	-- 3343
        b"010011000100_110001100000_000000100001_111110000000_000000000000_111000000000",	-- 3344
        b"010011110001_110001000000_000000100001_110001000001_011010100110_111010000000",	-- 3345
        b"010111001100_110000000000_000011101001_110011000010_011011101011_111000000000",	-- 3346
        b"110010000000_000000000000_000110100001_101110000000_000101111110_111000100000",	-- 3347
        b"010010001000_000000000000_000000100001_101110000000_000000011111_111000100000",	-- 3350
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3351
        b"110011000000_010100100000_000000100001_111110000000_000000000000_111010000000",	-- 3352
        b"110011001100_110000000000_000001101001_111011000010_001100010000_111000000000",	-- 3353
        b"010001101100_110000000000_000000100001_110001000001_011011001110_111000000000",	-- 3354
        b"010011001000_110010011000_000000100001_111011000001_001100010000_111000000000",	-- 3355
        b"110010000000_000000000000_000000100001_100001000001_011011110000_111000000000",	-- 3356
        b"010001101100_110101100000_000000100001_110011000001_100011111001_111000000000",	-- 3357
        b"010001101010_011000000000_000000100001_110001000001_011011001111_111000000000",	-- 3360
        b"110010000000_000000000000_000110100001_101110000000_000101111110_111000100000",	-- 3361
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3362
        b"011101101000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 3363
        b"110010000000_000000000000_000110100001_101110000000_000101110010_111000100000",	-- 3364
        b"010011111000_010100100000_000000100001_111110000000_000000000000_111000000000",	-- 3365
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3366
        b"010011110000_010100101000_000000100001_111010000001_000000000000_111000000000",	-- 3367
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3370
        b"010001101100_110010111000_000000100001_111011000001_001100010000_111000000000",	-- 3371
        b"010001101010_111101100000_000000100001_110011000001_100011111001_111000000000",	-- 3372
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3373
        b"110010000000_000000000000_000110100001_101110000000_000101111010_111000100000",	-- 3374
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3375
        b"110010000000_000000000000_000110100001_101110000000_000101111010_111000100000",	-- 3376
        b"010010000000_000101100000_000000100001_100011000001_100011111001_111010000000",	-- 3377
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3400
        b"110010000000_000000000000_000110100001_101110000000_000101111011_111000100000",	-- 3401
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3402
        b"110010000000_000000000000_000110100001_101110000000_000101111011_111000100000",	-- 3403
        b"010010000000_000101100000_000000100001_100011000001_100011111001_111010000000",	-- 3404
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3405
        b"110010000000_000000000000_000110100001_101110000000_000101111001_111000100000",	-- 3406
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3407
        b"110010000000_000000000000_000110100001_101110000000_000101111001_111000100000",	-- 3410
        b"010010000000_000101100000_000000100001_100011000001_100011111001_111010000000",	-- 3411
        b"110010000000_000000000000_101000100001_100001000001_011100001101_111000000000",	-- 3412
        b"110010000000_000000000000_100000100001_100001000001_011100001101_111000000000",	-- 3413
        b"110010000000_000000000000_000000100001_101011000001_001100010000_111000000000",	-- 3414
        b"110001101100_010000000001_111110100001_111110000000_000000000000_111000000000",	-- 3415
        b"110010001000_000000000000_000000100001_111010000001_000000000000_111010000000",	-- 3416
        b"010010001000_000101100000_000000100001_101110000000_000000011011_111000100000",	-- 3417
        b"010000010011_111101100010_000000100001_111110000000_000000000000_111000000000",	-- 3420
        b"010010001000_000001011000_000000100001_110001000001_011100011010_111000000000",	-- 3421
        b"110010000000_000000000000_000000100001_100001000001_011100011010_111000000000",	-- 3422
        b"110010000000_000000000000_000110100001_101110000000_000101110111_111000100000",	-- 3423
        b"100101101101_110101100000_010010100001_110001000001_011100011010_111000000000",	-- 3424
        b"010010000000_000101100000_000000100001_101110000000_000000000000_111010000000",	-- 3425
        b"110010000000_000000000000_000110100001_101110000000_000101110110_111000100000",	-- 3426
        b"010000110101_110001011000_000000100001_011110000000_000000000000_111000000000",	-- 3427
        b"010010000000_000101100000_000001001101_100011000011_100011111111_111010000000",	-- 3430
        b"010001101101_110101100010_000000100001_110011000001_100011111111_111000000000",	-- 3431
        b"100100110101_110101100000_010010100001_111110000000_000000000000_111000000000",	-- 3432
        b"010000110101_110001011000_000000100001_111010000001_000000000000_111000000000",	-- 3433
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3434
        b"110010000000_000000000000_000110100001_101110000000_000101110110_111000100000",	-- 3435
        b"110001101100_110000000000_000000100001_110001000001_100110110000_111010000000",	-- 3436
        b"110010000000_000000000000_000110100001_101110000000_000101110111_111000100000",	-- 3437
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3440
        b"110010000000_000000000000_000110100001_101110000000_000101110100_111000100000",	-- 3441
        b"010010000000_000101100000_000000100001_101110000000_000000000000_111010000000",	-- 3442
        b"100100110101_110101100000_010010100001_110011000001_100011111001_111000000000",	-- 3443
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3444
        b"110010000000_000000000000_000110100001_101110000000_000101110101_111000100000",	-- 3445
        b"000101101100_110100100010_000010100001_111110000000_000000000000_111000000000",	-- 3446
        b"000101101100_110100100010_000010100001_111110000000_000000000000_111010000000",	-- 3447
        b"110010000000_000000000000_000110100001_101110000000_000101110100_111000100000",	-- 3450
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3451
        b"011101101100_010100000001_111110100001_110001000001_100110110011_111000000000",	-- 3452
        b"110010000000_000000000000_000110100001_101110000000_000101101011_111000100000",	-- 3453
        b"110011000111_111100100000_011000100001_111011000001_001100010000_111010000000",	-- 3454
        b"110010000000_000000000000_000110100001_101110000000_000101101011_111000100000",	-- 3455
        b"010010000000_000101100000_000000100001_100011000001_100011111001_111010000000",	-- 3456
        b"110001101100_010000000000_000110100001_111110000000_000000000000_111000000000",	-- 3457
        b"010010000000_000101100000_000000100001_101110000000_000000000000_111001100000",	-- 3460
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111001100000",	-- 3461
        b"010010000000_010101101000_000000100001_100011000001_100011100010_111011100000",	-- 3462
        b"110011000111_110010100000_000000100001_011110000000_000000000000_111000000000",	-- 3463
        b"010010001000_000010000000_000000100001_101110000000_000010000000_111000100000",	-- 3464
        b"110001101010_110000000000_000111001001_110011000011_011100111001_111000000000",	-- 3465
        b"010010001000_000000000000_000000100001_101110000000_100010000000_111000100000",	-- 3466
        b"100100110000_010000000000_010010100001_111110000000_000000000000_111000000000",	-- 3467
        b"010010000000_010010001000_000000100001_101110000000_000000000000_111011100000",	-- 3470
        b"110001101010_010000000000_000000100001_110001000001_011101010100_111010000000",	-- 3471
        b"011001101010_110000000010_000110100001_111100000000_000000000101_111000000000",	-- 3472
        b"010010001000_000000010000_000000100001_111110000000_000000000000_111000000000",	-- 3473
        b"010010000000_000000001000_000000100001_100001000001_101000010000_111010000000",	-- 3474
        b"110001101000_000000000010_000110100001_111110000000_000000000000_111000000000",	-- 3475
        b"110010001000_000000000000_000000100001_111001000000_011100111101_111010000000",	-- 3476
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 3477
        b"010010001000_000000000000_000000100001_101110000000_000000011000_111000100000",	-- 3500
        b"010010001000_000000100000_000000100001_110001000001_011111001101_111000000000",	-- 3501
        b"110001101010_110000000010_000110100001_110001000001_001010001110_111000000000",	-- 3502
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3503
        b"010010001000_000000100000_000000100001_101110000000_000000010000_111000100000",	-- 3504
        b"010010000010_110001000000_000000100001_100001000001_011101001110_111011100000",	-- 3505
        b"110001101000_010000000000_000000100001_111110000000_000000000000_111010100000",	-- 3506
        b"010010001000_000000100000_000000100001_101110000000_000000001000_111000100000",	-- 3507
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 3510
        b"110000110010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3511
        b"010010000000_000000000000_000000100001_100001000001_011101001110_111010000000",	-- 3512
        b"110010000000_000000000000_000000100001_100001000001_011101010000_111000000000",	-- 3513
        b"110001101010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3514
        b"010010000000_000010000000_000000100001_100011000001_011101010100_111010000000",	-- 3515
        b"110000110000_110001000000_000110100001_111110000000_000000000000_111000000000",	-- 3516
        b"110001101000_010000000000_000000100001_111110000000_000000000000_111001100000",	-- 3517
        b"100100110000_010000000000_010010100001_111100000000_000000000011_111000000000",	-- 3520
        b"100100110000_010000000000_010010100001_111001000000_011101010001_111000000000",	-- 3521
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3522
        b"110001101000_010000000000_000000100001_111010000001_000000000000_111001100000",	-- 3523
        b"100101101010_010000100001_010010100001_111100000000_000000001000_111000000000",	-- 3524
        b"100101101000_110000100001_010010100001_111001000000_011101010101_111000000000",	-- 3525
        b"110011000111_110010100000_000000100001_011110000000_000000000000_111000000000",	-- 3526
        b"010010001000_000000000000_000000100001_101110000000_000000011000_111000100000",	-- 3527
        b"011001000010_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 3530
        b"110000111000_010000000000_000111001001_110011000010_011101011011_111000000000",	-- 3531
        b"110001101000_110000000000_000000100001_111010000001_000000000000_111001100000",	-- 3532
        b"010010001000_000000000000_000000100001_101110000000_000000000100_111000100000",	-- 3533
        b"110011110000_010000100000_000000100001_111010000001_000000000000_111001100000",	-- 3534
        b"110011000111_110010100000_000001101001_110011000011_011101101101_111000000000",	-- 3535
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 3536
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3537
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 3540
        b"010010000000_000000100000_000001101001_100011000010_011101101100_111010000000",	-- 3541
        b"010010001000_000000100000_000000100001_101110000000_000000000010_111000100000",	-- 3542
        b"110011000000_010000100000_000001101001_110011000011_011110010110_111000000000",	-- 3543
        b"110010000000_000000000000_000000100001_100001000001_001000000101_111000000000",	-- 3544
        b"110010000000_000000000000_000000100001_100001000001_011110101010_111000000000",	-- 3545
        b"110010000000_000000000000_000110100001_101110000000_000011000010_111000100000",	-- 3546
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3547
        b"110010000000_000000000000_000110100001_101110000000_000011000011_111000100000",	-- 3550
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 3551
        b"110010110000_010000100000_000001101001_110001000010_000111111100_111000000000",	-- 3552
        b"110010000000_000000000000_000000100001_100011000001_000110101110_111000000000",	-- 3553
        b"110011000100_111000000000_000001101001_110011000010_011110010110_111000000000",	-- 3554
        b"010010001000_000001100000_000000100001_101110000000_000000000100_111000100000",	-- 3555
        b"110001101010_010000000000_000001111101_110011000011_011101110100_111000000000",	-- 3556
        b"110000110010_110001100010_000110100001_111110000000_000000000000_111000000000",	-- 3557
        b"010010000000_000000000000_000001101001_100011000010_011110010110_111010000000",	-- 3560
        b"110010001000_000000000000_000000100001_110001000001_011110101010_111010000000",	-- 3561
        b"110010000000_000000000000_000000100001_100001000001_011110111000_111000000000",	-- 3562
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 3563
        b"010010001000_000000000000_000000100001_101110000000_000100000000_111000100000",	-- 3564
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3565
        b"110011000010_010000000000_000001101001_110011000010_011110010110_111000000000",	-- 3566
        b"010010001000_000000000000_000000100001_101110000000_011110010010_111000100000",	-- 3567
        b"110010000000_000000000000_000000100001_100001000001_101000001111_111000000000",	-- 3570
        b"110010000000_000000000000_000110100001_101110000000_000000011000_111000100000",	-- 3571
        b"010010000000_000000100000_000000100001_100001000001_011110011000_111010000000",	-- 3572
        b"100101101011_011000000001_010010100001_011110000000_000000000000_111000000000",	-- 3573
        b"100101101000_010000000001_010011011101_010011000011_011101111111_111000000000",	-- 3574
        b"110010000000_000000000000_000001011101_100011000011_011110000000_111000000000",	-- 3575
        b"110010000000_000000000000_000000100001_100011000001_011110000011_111000000000",	-- 3576
        b"010010000100_110100100000_000001011101_100011000010_011110000011_111011100000",	-- 3577
        b"100101101100_110100100000_010010100001_111100000000_000000000011_111000000000",	-- 3600
        b"100100110100_110100100000_010010100001_111001000000_011110000001_111000000000",	-- 3601
        b"010010000100_110100100000_000000100001_101110000000_000000000000_111011100000",	-- 3602
        b"010001101100_110000000000_000000100001_110001000001_011110101010_111000000000",	-- 3603
        b"110010000000_000000000000_000000101001_101011000011_011110001011_111000000000",	-- 3604
        b"110010000000_000000000000_000000100001_100001000001_011110111000_111000000000",	-- 3605
        b"010010001000_000001100000_000000100001_101110000000_000000000100_111000100000",	-- 3606
        b"110000110010_110001100000_000110100001_111110000000_000000000000_111000000000",	-- 3607
        b"010010000000_000011011000_000000100001_100001000001_100001000101_111010000000",	-- 3610
        b"110010000000_000000000000_000000100001_100001000001_011110011110_111000000000",	-- 3611
        b"110010000000_000000000000_000000101101_100001000010_011110101111_111000000000",	-- 3612
        b"110010000000_000000000000_000110100001_101110000000_000101010000_111000100000",	-- 3613
        b"110010001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 3614
        b"010010001000_000000000000_000000100001_110001000001_101000001111_111000000000",	-- 3615
        b"010001101110_010100011001_001100100001_111011000001_000011100010_111000000000",	-- 3616
        b"000101101101_111000000001_010010100001_111110000000_000000000000_111000000000",	-- 3617
        b"000101101000_010000000001_010010100001_111110000000_000000000000_111000000000",	-- 3620
        b"010011110000_010010000000_000000100001_110011000001_011110000101_111000000000",	-- 3621
        b"000101101101_111000000001_010010100001_111110000000_000000000000_111000000000",	-- 3622
        b"000101101000_010000000001_010010100001_111110000000_000000000000_111000000000",	-- 3623
        b"010011110000_010010000000_000000100001_110001000001_011110111000_111000000000",	-- 3624
        b"110010000000_000000000000_000000100001_100001000001_011110101111_111000000000",	-- 3625
        b"110010000000_000000000000_000000100001_100001000001_011110111111_111000000000",	-- 3626
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 3627
        b"110000110010_110001100010_000110100001_111110000000_000000000000_111000000000",	-- 3630
        b"010010000000_000011011000_000000100001_101110000000_000000000000_111010000000",	-- 3631
        b"010000010000_110011011010_000000100001_111110000000_000000000000_111010000000",	-- 3632
        b"110010010000_110011011000_000000100000_111110000000_000000000000_111000000000",	-- 3633
        b"000101101011_011011011001_010010100001_111110000000_000000000000_111000000000",	-- 3634
        b"000101101011_011011011001_010010100001_110011000001_100101111010_111000000000",	-- 3635
        b"110000110010_110001100000_000110100001_111110000000_000000000000_111000000000",	-- 3636
        b"010010000000_000011011000_000000100001_100001000001_100101111010_111010000000",	-- 3637
        b"110011000101_111100100000_000001101001_110011000011_001101100100_111000000000",	-- 3640
        b"010000000000_000011011010_001010100001_110001000001_100101111011_001001000000",	-- 3641
        b"110000110010_110001100000_000110100001_111110000000_000000000000_111000000000",	-- 3642
        b"010001101100_110011011000_000001101001_110011000010_001101100100_111010000000",	-- 3643
        b"010001101011_011011011010_001010100001_110001000001_100101111011_001001000000",	-- 3644
        b"110010000000_000000000000_000110100001_101110000000_000000011000_111000100000",	-- 3645
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 3646
        b"110010010000_010100100000_000001101001_110011000010_001101100100_111000000000",	-- 3647
        b"110000110010_110001100010_000110100001_111110000000_000000000000_111000000000",	-- 3650
        b"110011000111_111100100000_000000011100_111010000001_000000000000_111010000000",	-- 3651
        b"010010000010_110000100000_000000100001_101110000000_000000000000_111011100000",	-- 3652
        b"110001101000_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3653
        b"110001101000_010000000000_000000100001_111010000001_000000000000_111001100000",	-- 3654
        b"010010001000_000000000000_000000100001_101110000000_010000000000_111000100000",	-- 3655
        b"110001101010_110000000000_000110100001_110011000001_011110110001_111000000000",	-- 3656
        b"110001101010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3657
        b"010010001000_000000000000_000000100001_101110000000_000100000000_111000100000",	-- 3660
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3661
        b"010010010000_010010000000_000000100001_111010000001_000000000000_111010000000",	-- 3662
        b"010010001000_000000000000_000000100001_101110000000_000010000000_111000100000",	-- 3663
        b"110001101010_110000000000_000110100001_110011000001_011110111010_111000000000",	-- 3664
        b"010010001000_000000000000_000000100001_101110000000_000010000000_111000100000",	-- 3665
        b"110001101010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3666
        b"010010010000_010010000000_000000100001_110011000001_011010010101_111010000000",	-- 3667
        b"010010001000_000000000000_000000100001_101110000000_010000000000_111000100000",	-- 3670
        b"110001101010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 3671
        b"010011110000_010010000000_000000100001_110011000001_011010010101_111010000000",	-- 3672
        b"010010001000_000000000000_000000100001_101110000000_010000000000_111000100000",	-- 3673
        b"110001101010_110000000000_000110100001_110011000001_011110110111_111000000000",	-- 3674
        b"010001101101_111000100010_000000100001_110001000001_011111001001_111000000000",	-- 3675
        b"110011110000_010000100000_000000100001_111010000001_000000000000_111001100000",	-- 3676
        b"010001101101_111000100010_000000100001_110001000001_011111001001_111000000000",	-- 3677
        b"110010010000_110000000000_000000100001_111010000001_000000000000_111001100000",	-- 3700
        b"010010001000_000000100000_000000100001_101110000000_000000000100_111000100000",	-- 3701
        b"110010000000_000000000000_000000100001_100001000001_011111001001_111000000000",	-- 3702
        b"110011110000_010000100000_000000100001_111010000001_000000000000_111001100000",	-- 3703
        b"010010001000_000000100000_000000100001_101110000000_000000000100_111000100000",	-- 3704
        b"110010000000_000000000000_000000100001_100001000001_011111001001_111000000000",	-- 3705
        b"110010010000_110000000000_000000100001_111010000001_000000000000_111001100000",	-- 3706
        b"010010001000_000000000000_000000100001_101110000000_000000001000_111000100000",	-- 3707
        b"011101000010_110000000000_000000100001_100011000001_011111001011_111011100000",	-- 3710
        b"010010001000_000000000000_000000100001_101110000000_000000011000_111000100000",	-- 3711
        b"011101000010_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 3712
        b"110000111000_010000000000_000110100001_111110000000_000000000000_111000000000",	-- 3713
        b"010010000000_000000000000_000000100001_101010000001_000000000000_111001100000",	-- 3714
        b"011101000010_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 3715
        b"110000111000_010000000000_000110100001_111110000000_000000000000_111000000000",	-- 3716
        b"110001101000_110000000000_000000100001_111010000001_000000000000_111001100000",	-- 3717
        b"010010001000_000001100000_000000100001_101110000000_000000000110_111000100000",	-- 3720
        b"011110001010_110000000000_000000100001_100001000001_011111001011_111011100000",	-- 3721
        b"010010001000_000001000000_000000100001_101110000000_000011111111_111000100000",	-- 3722
        b"010011000000_010001000000_000000100001_110001000001_011111000111_111000000000",	-- 3723
        b"010010001000_000000100000_000000100001_101110000000_000000111000_111000100000",	-- 3724
        b"010011000000_110000000000_000001101001_010011000010_011111011001_111000000000",	-- 3725
        b"010010001000_000000100000_000000100001_101110000000_000100000000_111000100000",	-- 3726
        b"010011110000_110001000000_000000100001_111110000000_000000000000_111000000000",	-- 3727
        b"010010000000_010001001000_000000100001_101110000000_000000000000_111011100000",	-- 3730
        b"110011000111_110010100000_000001101001_110011000011_011111100000_111000000000",	-- 3731
        b"010010001000_000000100000_000000100001_101110000000_000001111111_111000100000",	-- 3732
        b"011111000001_010000100000_000000100001_101110000000_000000011100_111000100000",	-- 3733
        b"110010000000_000000000000_000110100001_101110000000_000011000000_111000100000",	-- 3734
        b"110000011000_110000000010_000001101001_110011000010_000111010010_111000000000",	-- 3735
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 3736
        b"110011000100_111000100000_000001101001_110011000010_000110010100_111000000000",	-- 3737
        b"110001101010_010000000000_000000100001_011110000000_000000000000_111000000000",	-- 3740
        b"110000110001_110010100000_000111011101_110011000011_011111101001_111000000000",	-- 3741
        b"110010000000_000000000000_000001101001_100011000010_011111100101_111010000000",	-- 3742
        b"010010001000_000000100000_000000100001_101110000000_000100010000_111000100000",	-- 3743
        b"010011110000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 3744
        b"010010000000_010001101000_000000100001_101110000000_000000000000_111011100000",	-- 3745
        b"110011000111_111001100000_000000100001_111110000000_000000000000_111010000000",	-- 3746
        b"110010000000_000000000000_000000100001_100001000001_011110110011_111000000000",	-- 3747
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 3750
        b"010010001000_000000000000_000000100001_101110000000_010000000000_111000100000",	-- 3751
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 3752
        b"110011000010_010000000000_000001101001_110011000010_100000000100_111000000000",	-- 3753
        b"010010001000_000000000000_000000100001_101110000000_100000001000_111000100000",	-- 3754
        b"110010000000_000000000000_000000100001_100001000001_101000001111_111000000000",	-- 3755
        b"110010000000_000000000000_000110100001_101110000000_000000011000_111000100000",	-- 3756
        b"010010000000_000000100000_000000100001_100001000001_011110011000_111010000000",	-- 3757
        b"010010001000_000000000000_000000100001_101110000000_000111111111_111000100000",	-- 3760
        b"100101101011_011000100001_010010100001_011110000000_000000000000_111000000000",	-- 3761
        b"100101101000_110000100001_010011011101_010011000011_011111110101_111000000000",	-- 3762
        b"110010000000_000000000000_000001011101_100011000011_011111110111_111000000000",	-- 3763
        b"110010000000_000000000000_000000100001_100011000001_011111111011_111000000000",	-- 3764
        b"010010000001_010001000000_000000100001_101110000000_000000000000_111011100000",	-- 3765
        b"010010000000_010000000000_000001011101_100011000010_011111111011_111011100000",	-- 3766
        b"100101101001_010001000000_010010100001_111110000000_000000000000_111000000000",	-- 3767
        b"100101101000_010000000000_010010100001_111100000000_000000000011_111000000000",	-- 3770
        b"100100110001_010001000000_010010100001_111110000000_000000000000_111000000000",	-- 3771
        b"100100110000_010000000000_010010100001_111001000000_011111111001_111000000000",	-- 3772
        b"010010010000_010100100000_000000100001_111110000000_000000000000_111000000000",	-- 3773
        b"010011110001_010100100000_000000100001_110001000001_100111000100_111000000000",	-- 3774
        b"110010000000_000000000000_000000101001_100011000011_100000000100_111000000000",	-- 3775
        b"110010000000_000000000000_000000100001_100001000001_011110110011_111000000000",	-- 3776
        b"010010001000_000001100000_000000100001_101110000000_000000000110_111000100000",	-- 3777
        b"110000110010_110001100000_000110100001_111110000000_000000000000_111000000000",	-- 4000
        b"010010000000_000011011000_000000100001_100001000001_100001000101_111010000000",	-- 4001
        b"110010000000_000000000000_000000100001_100001000001_011110011110_111000000000",	-- 4002
        b"110010000000_000000000000_000000101101_100001000010_011110101101_111000000000",	-- 4003
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 4004
        b"000101101101_111000000001_010010100001_111100000000_000000000001_111000000000",	-- 4005
        b"000101101000_010000000001_010010100001_111001000000_100000000110_111000000000",	-- 4006
        b"010011110000_010010000000_000000100001_110011000001_011111111110_111000000000",	-- 4007
        b"000101101101_111000000001_010010100001_110100000001_000000000001_111000000000",	-- 4010
        b"000101101000_010000000001_010010100001_111000000000_000000000000_111000000000",	-- 4011
        b"010011110000_010010000000_000000100001_110001000001_011110110011_111000000000",	-- 4012
        b"110010000000_000000000000_000000100001_100011000001_011110001011_111000000000",	-- 4013
        b"110010000000_000000000000_000000100001_100001000001_011111000111_111000000000",	-- 4014
        b"010010001000_000000100000_000000100001_101110000000_000011000000_111000100000",	-- 4015
        b"010011000000_110000000000_000000100001_110001000001_100000010111_111000000000",	-- 4016
        b"011011000000_110010000000_000000100001_100001000001_011000011001_111000000000",	-- 4017
        b"110010111000_010000000000_000001101001_110011000010_100000010101_111000000000",	-- 4020
        b"010010010000_110010000000_000000100001_111110000000_000000000000_111000000000",	-- 4021
        b"010010001000_000000110000_000000100001_101110000000_100000000000_111000100000",	-- 4022
        b"100100110000_110000110000_010010100001_111110000000_000000000000_111000000000",	-- 4023
        b"110011110000_110010000000_000000100001_111110000000_000000000000_111010000000",	-- 4024
        b"110010000000_000000000000_000000100001_101011000001_011110001011_111000000000",	-- 4025
        b"010010000000_010000000000_000000100001_101010000001_000000000000_111011100000",	-- 4026
        b"010010000000_110000100000_000000100001_101010000001_000000000000_111011100000",	-- 4027
        b"110010000000_000000000000_000000100001_100001011110_011000111010_111000000000",	-- 4030
        b"110010000000_000000000000_000000100001_100110000001_100100000000_111000000000",	-- 4031
        b"110011000101_010101100000_011001101001_111011000011_001100010000_111000000000",	-- 4032
        b"010001101011_110011110010_000000100001_111011000001_001100010000_111000000000",	-- 4033
        b"110011000101_010101100000_011001101001_110011000010_001100010000_111000000000",	-- 4034
        b"010001101011_110011110010_000000100001_111011000001_001100010000_111000000000",	-- 4035
        b"010010000000_000101100000_000000100001_100011000001_100000011111_111010000000",	-- 4036
        b"110010000000_000000000000_000000100001_100001000001_100000100010_111000000000",	-- 4037
        b"110010000000_000000000000_011000101101_101011000011_001100010000_111000000000",	-- 4040
        b"110010000000_000000000000_000000100001_101011000001_100111100101_111000000000",	-- 4041
        b"010011000110_111100000000_000000011110_110001000001_001101100101_111000000000",	-- 4042
        b"010001101100_010011011000_001011011101_110011000010_100000100111_100001000000",	-- 4043
        b"010001101101_110101100000_001010100001_011110000000_000000000000_101001000000",	-- 4044
        b"110010000000_000000000000_000000011100_101010110001_000000000000_000000000000",	-- 4045
        b"110010000000_000000000000_000000011110_101010000001_000000000000_111000000000",	-- 4046
        b"110000100100_010000000010_000001111101_011010000010_000000000000_111000000000",	-- 4047
        b"010010000000_000001000000_000001001001_100011000010_100001010100_111010000000",	-- 4050
        b"010001101101_110010000000_000000011100_111110000000_000000000000_111010000000",	-- 4051
        b"011011000000_110100000000_000001101001_110011000010_100000110001_111000000000",	-- 4052
        b"010010001000_000000100000_000000100001_101110000000_000000000101_111000100000",	-- 4053
        b"110000011000_110000000010_000000100001_011110000000_000000000000_111000000000",	-- 4054
        b"010010010000_010010100000_000001101001_110011000010_100001010001_111000000000",	-- 4055
        b"011000111111_111000000000_000001101001_110011000010_100000110000_111000000000",	-- 4056
        b"011000111111_111000000000_000001101001_111010000011_000000000000_111000000000",	-- 4057
        b"110010000000_000000000000_000000100001_100011000001_011101000000_111000000000",	-- 4060
        b"010010001000_000000000000_000000100001_101110000000_100000000000_111000100000",	-- 4061
        b"100101101000_010000000001_010010100001_111110000000_000000000000_111000000000",	-- 4062
        b"110011000000_010101100000_000001101001_110011000011_011100110011_111000000000",	-- 4063
        b"110010000000_000000000000_000110100001_101110000000_000101100001_111000100000",	-- 4064
        b"010010110010_010001000000_000000100001_111110000000_000000000000_111010000000",	-- 4065
        b"110010000000_000001000000_000000100001_100001101100_100001000000_111000000000",	-- 4066
        b"110010000000_000000000000_000110100001_101110000000_000001000111_111000100000",	-- 4067
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 4070
        b"110011000000_010001000000_000001101001_110001000011_100000111100_111000000000",	-- 4071
        b"110010000000_000000000000_000000100001_100001000001_011101010100_111000000000",	-- 4072
        b"110010000000_000000000000_000000011100_100011000001_011010010101_111000000000",	-- 4073
        b"010010001000_000001100000_000000100001_101110000000_000000000110_111000100000",	-- 4074
        b"110000110010_110001100000_000110011110_111110000000_000000000000_111000000000",	-- 4075
        b"110011000000_010010000000_000001101001_110011000011_100001001010_111000000000",	-- 4076
        b"110010000000_000000000000_000000100001_100011000001_100001000101_111000000000",	-- 4077
        b"010010001000_000000000000_000000100001_101110000000_000100000000_111000100000",	-- 4100
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 4101
        b"010010001000_000001100000_000000100001_101110000000_000000000100_111000100000",	-- 4102
        b"110000110010_110001100000_000110011110_111110000000_000000000000_111000000000",	-- 4103
        b"110011000000_010010000000_000001101001_110011000011_100001001101_111000000000",	-- 4104
        b"110000110010_110001100010_000110100001_111110000000_000000000000_111000000000",	-- 4105
        b"010010000000_000100100000_000000100001_100001000001_011100001110_111010000000",	-- 4106
        b"010001101011_011011011010_000000100001_110001000001_100111000100_111000000000",	-- 4107
        b"110010000000_000000000000_000110100001_101110000000_000101100001_111000100000",	-- 4110
        b"010010000000_000001000000_000000100001_101010000001_000000000000_111010000000",	-- 4111
        b"010010000000_000011011000_000001101001_100001000011_011110100100_111010000000",	-- 4112
        b"110010000000_000000000000_000000101101_100001000010_011110101101_111000000000",	-- 4113
        b"110010000000_000000000000_000000100001_100011000001_100001001111_111000000000",	-- 4114
        b"010010000000_000011011000_000001101001_100001000011_011110100100_111010000000",	-- 4115
        b"110010000000_000000000000_000000101101_100001000010_011110101111_111000000000",	-- 4116
        b"110010000000_000000000000_000110100001_101110000000_000101100001_111000100000",	-- 4117
        b"010010000000_000001000000_000000100001_101010000001_000000000000_111010000000",	-- 4120
        b"110010000000_000000000000_000000100001_100001000001_011110111101_111000000000",	-- 4121
        b"110001101010_110000000000_000110100001_111110000000_000000000000_111000000000",	-- 4122
        b"010010000000_000010000000_000000100001_100011000001_011110111011_111010000000",	-- 4123
        b"110001101101_110000000000_000000011100_111010000001_000000000000_111010000000",	-- 4124
        b"010011110101_010101100000_000000100001_111011000001_100000011111_111000000000",	-- 4125
        b"010010010101_010101100000_000000100001_111011000001_100000011111_111000000000",	-- 4126
        b"110010000000_000000000000_011000100001_101011110111_001100010000_111000000000",	-- 4127
        b"010010001000_000000000001_110000100001_101110000000_000110000000_111000100000",	-- 4130
        b"010010000000_010011011000_011000100001_101011100001_001100010000_111011100000",	-- 4131
        b"010011000000_011011011000_000001101001_111011000010_001100010000_111000000000",	-- 4132
        b"110010000000_000000000000_000000100001_100100000001_000000001000_111000000000",	-- 4133
        b"100101101011_011011011001_010010100001_111000000000_000000000000_111000000000",	-- 4134
        b"010010001000_000000000000_000000100001_101110000000_000100010000_111000100000",	-- 4135
        b"010000110000_010011011000_000000100001_110001000001_100001100000_111000000000",	-- 4136
        b"110010000000_000000000000_000000100001_100011000001_001100011101_111000000000",	-- 4137
        b"110010000000_000000000000_000000100001_100011011111_100001100010_111000000000",	-- 4140
        b"010000110010_011011011000_001010100001_110011000001_100101111011_001001000000",	-- 4141
        b"010000110001_111011011000_001010100001_110011000001_100101111011_001001000000",	-- 4142
        b"010010001000_000000000001_111000100001_101110000000_100000000010_111000100000",	-- 4143
        b"010010000000_010000000000_000000100001_100011000001_100001101001_111011100000",	-- 4144
        b"010010001000_000000000001_111000100001_101110000000_000010000000_111000100000",	-- 4145
        b"010010000000_010000000000_000000100001_100011000001_100001101011_111011100000",	-- 4146
        b"010010001000_000000000001_111000100001_101110000000_000100000000_111000100000",	-- 4147
        b"010010000000_010000000000_000000100001_100011000001_100001101011_111011100000",	-- 4150
        b"100100110000_010000000000_010010100001_111100000000_000000000001_111000000000",	-- 4151
        b"100100110000_010000000000_010010100001_111001000000_100001101010_111000000000",	-- 4152
        b"010011110000_010000011000_000000100001_111010000001_000000000000_111000000000",	-- 4153
        b"010000110111_111011111000_101100100001_011011111100_100010010110_000000000000",	-- 4154
        b"110001101100_011000000001_001101001001_111010000011_000000000000_000000000000",	-- 4155
        b"110010000000_000000000000_000110100001_101110000000_000101011101_111000100000",	-- 4156
        b"110011000111_111000100000_000000100001_111110000000_000000000000_111010000000",	-- 4157
        b"110010000000_000000000000_000110100001_101110000000_000101011110_111000100000",	-- 4160
        b"110011000111_111001000000_000000100001_111110000000_000000000000_111010000000",	-- 4161
        b"010010001000_000011111000_000000100001_101110000000_000000011011_111000100000",	-- 4162
        b"110010000000_000000000000_000110100001_101110000000_000101110111_111000100000",	-- 4163
        b"010010001000_000000100000_000000100001_101110000000_111110100000_111000100000",	-- 4164
        b"011101101000_110000100000_000000100001_101110000000_000000000000_111010000000",	-- 4165
        b"011000111000_110000000000_000001101101_110011000011_100001111100_111010000000",	-- 4166
        b"000110001000_000000100000_001010100001_101110000000_000000000000_111000100000",	-- 4167
        b"110000111000_110000000000_000000100001_111110000000_000000000000_111010000000",	-- 4170
        b"110010000000_000000000000_000110100001_101110000000_000101110110_111000100000",	-- 4171
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 4172
        b"110001101000_110000000010_000000100001_111110000000_000000000000_111010000000",	-- 4173
        b"110010000000_000000000000_000110100001_101110000000_000101110100_111000100000",	-- 4174
        b"010010000000_000000100000_000000100001_001110000000_000000000000_111010000000",	-- 4175
        b"110010000000_000000000000_000110100001_101110000000_000101110101_111000100000",	-- 4176
        b"011101101000_110000100000_000001001001_100011000010_100010010001_111010000000",	-- 4177
        b"110000110111_111000100000_000001101001_110011000011_100010010001_111010000000",	-- 4200
        b"110011001111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 4201
        b"110010000000_000000000000_000110100001_101110000000_000101101110_111000100000",	-- 4202
        b"010010001000_000000100000_000000100001_101110000000_000000100000_111000100000",	-- 4203
        b"011101101000_010000100000_000000100001_101110000000_000000000000_111010000000",	-- 4204
        b"010011111000_110000100000_000000100001_111110000000_000000000000_111010000000",	-- 4205
        b"010010000000_110001000000_000000100001_101110000000_000000000000_111011100000",	-- 4206
        b"110011000000_110001000000_000000100001_011110000000_000000000000_111000000000",	-- 4207
        b"010010001000_000001000000_000000100001_101110000000_000000000111_111000100000",	-- 4210
        b"010011000000_110001000000_000001001001_010011000010_100010010001_111000000000",	-- 4211
        b"010010001000_000000100000_000000100001_101110000000_000001011100_111000100000",	-- 4212
        b"110000110000_110001000000_000111001001_110011000010_100010010001_111000000000",	-- 4213
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 4214
        b"110010000000_000000000000_000110100001_101110000000_000101110011_111000100000",	-- 4215
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 4216
        b"110001101001_010000000000_000000100001_111110000000_000000000000_111010000000",	-- 4217
        b"110011110000_110001000000_000000100001_111110000000_000000000000_111100000000",	-- 4220
        b"110010000000_000000000000_000110100001_101110000000_000101011101_111000100000",	-- 4221
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 4222
        b"110010000000_000000000000_000110100001_101110000000_000101011110_111000100000",	-- 4223
        b"010010000000_000001000000_000000100001_101110000000_000000000000_111010000000",	-- 4224
        b"010001101011_011011011000_001010100001_111010000001_000000000000_001001000000",	-- 4225
        b"010001101011_111011111010_000000100001_111011100011_100010011000_111000000000",	-- 4226
        b"010000110111_111011110000_000000100001_111101000001_000000000000_111000000000",	-- 4227
        b"010001101100_011110000000_011000100001_111101000001_000000000000_111000000000",	-- 4230
        b"010010000000_000100011000_110100100001_101101000001_000000000000_111000000000",	-- 4231
        b"010010001000_000010100000_000000100001_101101000001_000000000111_111000100000",	-- 4232
        b"010011000010_110110000000_000000100001_111110000000_000000000000_111000000000",	-- 4233
        b"110010110010_110110000000_000001101001_110011000010_100010011100_111000000000",	-- 4234
        b"010011000010_110100011000_000000100001_111101000001_000000000000_111000000000",	-- 4235
        b"110010000000_000000000000_000000100001_100001100110_010100010100_111000000000",	-- 4236
        b"110010110010_110100011000_000001101001_110011000011_100010110010_111000000000",	-- 4237
        b"110010000000_000000000000_000110100001_101110000000_000101010000_111000100000",	-- 4240
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 4241
        b"010001101000_010000000000_000001101001_110011000011_100010100010_111000000000",	-- 4242
        b"110000001000_000000000000_000000100001_111110000000_000000000000_111010000000",	-- 4243
        b"010001101000_001000000000_000000100001_111101000001_000000000000_111000000000",	-- 4244
        b"010010001000_000000100000_000000100001_101110000000_000001000000_111000100000",	-- 4245
        b"110011000000_010000100000_000001101001_110011000011_100010100110_111000000000",	-- 4246
        b"010011000000_010010100000_000000100001_111110000000_000000000000_111000000000",	-- 4247
        b"010010000010_110010101000_000000100001_101110000000_000000000000_111011100000",	-- 4250
        b"100100110010_110010110000_010010100001_111110000000_000000000000_111000000000",	-- 4251
        b"011100110010_110010110000_000000100001_101110000000_000010000000_111000100000",	-- 4252
        b"010000111010_110010110000_000110100001_111110000000_000000000000_111000000000",	-- 4253
        b"010010000000_000010000000_000000100001_101110000000_000000000000_111010000000",	-- 4254
        b"010010001000_000000100000_000000100001_101110000000_000000001000_111000100000",	-- 4255
        b"110011000000_010000100000_000001101001_111011000011_011101011101_111000000000",	-- 4256
        b"010010001000_000000100000_000000100001_101110000000_000000010000_111000100000",	-- 4257
        b"110011000000_010000100000_000001101001_111011000010_011111010000_111000000000",	-- 4260
        b"110010000000_000000000000_000000100001_101011000001_100000001100_111000000000",	-- 4261
        b"010010001000_000000000000_000000100001_101110000000_000001100100_111000100000",	-- 4262
        b"110000100000_010100011000_000110100001_110001000001_001010001110_111000000000",	-- 4263
        b"110010000000_000000000000_000110100001_101110000000_000101101111_111000100000",	-- 4264
        b"011101101000_010000000000_000000100001_101110000000_000000000000_111010000000",	-- 4265
        b"110011111000_010000000000_000000100001_111110000000_000000000000_111010000000",	-- 4266
        b"010010001000_000100000000_000000100001_101110000000_000000110000_111000100000",	-- 4267
        b"011000100100_010100011000_000110100001_101110000000_000000010111_111000100000",	-- 4270
        b"011100011100_011010000010_000000100001_100011100100_100010111011_111010000000",	-- 4271
        b"010001110111_110010000000_000000100001_111110000000_000000000000_111000000000",	-- 4272
        b"010010001000_000000000000_000000100001_101110000000_100011001111_111000100000",	-- 4273
        b"110010000000_000000000000_000000100001_100001000001_101000001111_111000000000",	-- 4274
        b"010000111001_111011011000_001010100001_110001000001_100101111011_001001000000",	-- 4275
        b"010001101100_110100000000_000000100001_011110000000_000000000000_111000000000",	-- 4276
        b"110010010010_010100100000_000001001001_010011000010_100011001111_111000000000",	-- 4277
        b"010001101000_011100100000_000000100001_111110000000_000000000000_111000000000",	-- 4300
        b"000101101100_111000000001_010010100001_110001000001_100011010001_111000000000",	-- 4301
        b"000101101000_010000000001_010010100001_110001000001_100011010001_111000000000",	-- 4302
        b"110010000000_000000000000_000000100001_100001011110_100001101011_111000000000",	-- 4303
        b"010011000110_111011100000_100001001001_110011000010_100011010010_111000000000",	-- 4304
        b"010010001000_000000000000_000000100001_101110000000_000010110100_111000100000",	-- 4305
        b"010010000000_010000000000_000000100001_100001000001_011011001111_111011100000",	-- 4306
        b"110011000111_110011100000_000000100001_010011100100_100011001111_111000000000",	-- 4307
        b"010010110000_010100000000_000001001001_110011000011_100011001111_111000000000",	-- 4310
        b"110011000111_110100000000_000001101001_110011000011_100011001111_111000000000",	-- 4311
        b"110010000000_000000000000_000110100001_101110000000_000001100101_111000100000",	-- 4312
        b"010010000000_000000000000_000000100001_100001000001_100011010001_111010000000",	-- 4313
        b"010001101011_110100110000_000000100001_110001000001_100111001001_111000000000",	-- 4314
        b"010010001000_000000000000_000000100001_110001000001_101000001111_111000000000",	-- 4315
        b"010001101100_010011110010_011000100001_111011000001_001100010000_111000000000",	-- 4316
        b"010010001000_000000000000_000000100001_101110000000_000001000001_111000100000",	-- 4317
        b"110010000000_000000000000_000000100001_101011000001_001001110110_111000000000",	-- 4320
        b"010010010000_010000011000_000000100001_111010000001_000000000000_111000000000",	-- 4321
        b"010001101000_010010000000_000000100001_110001000001_100111001001_111000000000",	-- 4322
        b"010001101011_110100100000_010000100001_110001000001_100111001000_111000000000",	-- 4323
        b"011101101100_010100000011_111110100001_110001000001_100110110011_111000000000",	-- 4324
        b"000101101100_111000000001_010010100001_110001000001_100011011011_111000000000",	-- 4325
        b"010010010010_010100100000_000000100001_111110000000_000000000000_111000000000",	-- 4326
        b"010011000010_010000011000_000000100001_111110000000_000000000000_111000000000",	-- 4327
        b"010011110100_110000011000_000000100001_110001000001_100110110000_111000000000",	-- 4330
        b"010010001000_000000000000_000000100001_110001000001_101000001111_111000000000",	-- 4331
        b"010001101100_110011100000_011000100001_111011000001_001100010000_111000000000",	-- 4332
        b"010010010000_010100100000_000000100001_111010000001_000000000000_111000000000",	-- 4333
        b"010001101101_110100100000_000000100001_110011100111_100011011111_111000000000",	-- 4334
        b"110010000000_000000000000_000000100001_100001000001_010100001011_111000000000",	-- 4335
        b"110010000000_000000000000_000000100001_100011000001_100011100000_111000000000",	-- 4336
        b"011111000110_111100000001_111110010110_110001000001_100111001010_111000000000",	-- 4337
        b"110010000000_000000000000_101110100001_101110000000_000000010000_111000000000",	-- 4340
        b"110011000111_111001011000_000000100001_110011000001_100011100010_111010000000",	-- 4341
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 4342
        b"110011000111_111101100000_011000100001_111011110111_001100010000_111010000000",	-- 4343
        b"110010000000_000000000000_000000100001_101011000001_100001011000_111000000000",	-- 4344
        b"110011000111_111101100000_101110100001_111110000000_000000010000_111010000000",	-- 4345
        b"110011000111_111001011000_011000100001_110011110111_001100010000_111010000000",	-- 4346
        b"110010000000_000000000000_000000100001_101011000001_100001011000_111000000000",	-- 4347
        b"110011000111_111101000000_011000100001_111011110111_001100010000_111010000000",	-- 4350
        b"110010000000_000000000000_000000100001_101011000001_100001011000_111000000000",	-- 4351
        b"010001101011_011011011000_001010100001_110011010011_100011101101_010001000000",	-- 4352
        b"010001101101_110101100000_001010100001_010011000110_100011111000_101001000000",	-- 4353
        b"010001101101_110100100000_000000100001_110011110001_100001010111_000010000000",	-- 4354
        b"110010000000_000000000000_000000100001_100011000110_100011111001_111000000000",	-- 4355
        b"110011000111_111101100000_000000100001_110011000001_100011111001_111010000000",	-- 4356
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 4357
        b"110011000111_111101100000_000000100001_110011000001_100011111001_111010000000",	-- 4360
        b"110011000111_111101100000_000000100001_111110000000_000000000000_111010000000",	-- 4361
        b"010001101101_010101100000_000000100001_111110000000_000000000000_111000000000",	-- 4362
        b"010001101011_011011011000_001010100001_110011010010_100011110111_010001000000",	-- 4363
        b"110001101011_011000000000_100110100001_110011100110_100011111001_111000000000",	-- 4364
        b"110011000111_111101100000_011000100001_111011110111_001100010000_111010000000",	-- 4365
        b"110010000000_000000000000_000000100001_100011000001_100001011000_111000000000",	-- 4366
        b"010001101101_110101100000_001010100001_011110000000_000000000000_101001000000",	-- 4367
        b"110010000000_000000000000_011000100001_100011110001_100001010111_000000000000",	-- 4370
        b"010001101101_110100100000_000000100001_110011100110_100011111101_111000000000",	-- 4371
        b"011111000110_111100000001_111110010110_110001000001_100111001010_111000000000",	-- 4372
        b"110010000000_000000000000_011000100001_100011110111_001100010000_111000000000",	-- 4373
        b"110010000000_000000000000_000000100001_100011000001_100001011000_111000000000",	-- 4374
        b"110010000000_000000000000_000000100001_100001000001_010100001011_111000000000",	-- 4375
        b"110010000000_000000000000_000000100001_101011000001_100001010111_111000000000",	-- 4376
        b"010001101101_110100100000_000000100001_110011100110_100100000100_111000000000",	-- 4377
        b"011111000110_111100000001_111110010110_110001000001_100111001010_111000000000",	-- 4400
        b"010001101001_011100100000_000000100001_110001000001_100111001000_111000000000",	-- 4401
        b"110010000000_000000000000_011000100001_100011110111_001100010000_111000000000",	-- 4402
        b"110010000000_000000000000_000000100001_100011000001_100001011000_111000000000",	-- 4403
        b"010010001000_000110010000_000000100001_101110000000_000010000000_111000100000",	-- 4404
        b"110010000000_000000000000_000000100001_100001000001_010100011010_111000000000",	-- 4405
        b"011111000110_111100000001_111110010110_110001000001_100111001010_111000000000",	-- 4406
        b"010001101001_011100100000_000000100001_110001000001_100111001000_111000000000",	-- 4407
        b"110010000000_000000000000_000000100001_100001000001_010100010100_111000000000",	-- 4410
        b"110010000000_000000000000_000000100001_101011000001_100001010111_111000000000",	-- 4411
        b"110010000000_000000000000_101110100001_101110000000_000000000000_111000000000",	-- 4412
        b"110011000111_111101100000_101110100001_111110000000_000000010000_111010000000",	-- 4413
        b"110011000111_111001011000_101110100001_111110000000_000000100000_111010000000",	-- 4414
        b"110011000111_111101000000_101110100001_111110000000_000000110000_111010000000",	-- 4415
        b"110011000111_111000111000_011000100001_111011110111_001100010000_111010000000",	-- 4416
        b"110010000000_000000000000_000000100001_101011000001_100001011000_111000000000",	-- 4417
        b"010010001000_000000000000_000000100001_101100000000_000111111111_111000100000",	-- 4420
        b"010001101000_010000000010_000110100001_111110000000_000000000000_111000000000",	-- 4421
        b"110010001000_000000000000_000000100001_111001000000_100100010001_111010000000",	-- 4422
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 4423
        b"110010000000_000000000000_000110010110_101110000000_000100100001_111000100000",	-- 4424
        b"110011000111_111100100000_000000100001_110011000001_100100010110_111010000000",	-- 4425
        b"110010000000_000000000000_000000100001_100011100101_100101010110_111000000000",	-- 4426
        b"010010000100_010011011000_000000100001_101011010101_100111101001_111011100000",	-- 4427
        b"010011000110_110011011000_000000100001_110011011111_100100011010_111000000000",	-- 4430
        b"010000110010_011011011000_000000100001_110011000001_100100011011_111000000000",	-- 4431
        b"010000110001_111011011000_000000100001_111110000000_000000000000_111000000000",	-- 4432
        b"010010001000_000000000000_000000100001_101110000000_000101100000_111000100000",	-- 4433
        b"010001101100_111001000000_000000010000_111110000000_000000000000_111000000000",	-- 4434
        b"011100110000_010011011000_001010100001_110001000001_100100110011_001001000000",	-- 4435
        b"010001101100_110000100000_000000100001_110001000001_100101000111_111000000000",	-- 4436
        b"100101101100_010000000000_010010100001_110100000001_000000000011_111000000000",	-- 4437
        b"100100110000_010000000000_010010100001_111000000000_000000000000_111000000000",	-- 4440
        b"010010000000_010011011000_000000100001_101110000000_000000000000_111011100000",	-- 4441
        b"010011000111_010011011000_000000100001_111110000000_000000000000_111000000000",	-- 4442
        b"010000110001_110011011000_001010100001_110001000001_100100110011_001001000000",	-- 4443
        b"010001101100_110000100000_000000010010_110001000001_100101000111_111000000000",	-- 4444
        b"010010001000_000000000000_000000100001_101110000000_000000000001_111000100000",	-- 4445
        b"110011000100_110000000000_000000100001_011110000000_000000000000_111000000000",	-- 4446
        b"011000110001_010001000000_000001001001_100011000010_100100101001_111000000000",	-- 4447
        b"010011111001_010001000000_000000100001_111110000000_000000000000_111000000000",	-- 4450
        b"011011110001_010001100000_000110100001_101110000000_000001000010_111000100000",	-- 4451
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 4452
        b"010011111000_010100100000_000000100001_110001011110_101000001010_111000000000",	-- 4453
        b"110001101100_010000000001_111110100001_111110000000_000000000000_111000000000",	-- 4454
        b"000110001000_000000100000_001010100001_101110000000_001111111110_111000100000",	-- 4455
        b"000101101000_110000100001_010010100001_111110000000_000000000000_111000000000",	-- 4456
        b"110011000100_110000100000_000001101001_110011000011_100111101101_111000000000",	-- 4457
        b"010001101100_110000000000_000000110101_111010000011_000000000000_111010000000",	-- 4460
        b"110010000000_000000000000_000110100001_101110000000_000100100001_111000100000",	-- 4461
        b"010010000000_000100100000_000000100001_101010000001_000000000000_111010000000",	-- 4462
        b"110010000000_000000000000_000000100001_100001000001_100101111011_000000000000",	-- 4463
        b"010011000100_110001000000_000000100001_111110000000_000000000000_111000000000",	-- 4464
        b"100101101100_110001100000_010010100001_011110000000_000000000000_111000000000",	-- 4465
        b"100101101001_110001100000_010011011101_010011000010_100111100100_111000000000",	-- 4466
        b"100101101001_110001100000_010011011101_010011000011_100101000000_111000000000",	-- 4467
        b"011010010111_110100100000_000001011101_100011000011_100100111101_111000000000",	-- 4470
        b"010010000100_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 4471
        b"010011000111_010000000000_000000100001_110001000001_100100111101_111000000000",	-- 4472
        b"010001101001_110011011000_000000100001_111110000000_000000000000_111000000000",	-- 4473
        b"010000110000_010011011000_001010100001_110011000001_100100110011_001001000000",	-- 4474
        b"011100111010_111011011000_001010100001_111110000000_000000000000_001001000000",	-- 4475
        b"110010000000_000000000000_000000100001_100001000001_100101111011_111000000000",	-- 4476
        b"100101101100_110001100000_010010000011_010001000001_100101000101_111000000000",	-- 4477
        b"100100110001_110001100000_010011011101_110011000011_100111100100_111000000000",	-- 4500
        b"010010000110_110000000000_000000100001_101110000000_000000000000_111011100000",	-- 4501
        b"110011000100_110000000000_000000100001_011110000000_000000000000_111000000000",	-- 4502
        b"010001101100_010001101000_000001001001_110011000011_100111100100_111000000000",	-- 4503
        b"100100110001_110001100000_010010100001_111110000000_000000000000_111000000000",	-- 4504
        b"100100110001_110001100000_010010100001_111110000000_000000000000_111000000000",	-- 4505
        b"110010000000_000000000000_000000100001_101010000001_000000000000_111000000000",	-- 4506
        b"110010000000_000000000000_000110100001_101110000000_000101111001_111000100000",	-- 4507
        b"010010001000_000011011000_000000100001_101110000000_111111111111_111000100000",	-- 4510
        b"100111000111_111011011000_011010100001_111110000000_000000000000_111000000000",	-- 4511
        b"011111000100_110011011000_000000100001_101110000000_000000000000_111010000000",	-- 4512
        b"010000111011_011011011000_001010100001_110001000001_100101111011_001001000000",	-- 4513
        b"110010000000_000000000000_000110100001_101110000000_000101111010_111000100000",	-- 4514
        b"110010010110_111100100000_000000100001_011110000000_000000000000_111000000000",	-- 4515
        b"011101101100_110100100000_000001001001_100011000010_100111100010_111010000000",	-- 4516
        b"011011001100_110000000000_000110100001_101110000000_000101111011_111000100000",	-- 4517
        b"010010000000_000100100000_000000100001_101110000000_000000000000_111010000000",	-- 4520
        b"011111111100_110100100000_000000110101_110011000011_100101010101_111000000000",	-- 4521
        b"110001101001_010000000000_000000101001_010011000011_100101010101_111000000000",	-- 4522
        b"010010001000_000100100000_000000100001_101110000000_000000000001_111000100000",	-- 4523
        b"010011111100_110100100000_000001001001_110011000010_100111100100_111000000000",	-- 4524
        b"010001101011_011011011000_001010100001_110011000001_100111000100_010001000000",	-- 4525
        b"110011000111_110100000000_000001101001_111011000011_100111101001_111000000000",	-- 4526
        b"011010010111_010100000000_000000100001_101110000000_000000000000_111000000000",	-- 4527
        b"010011001111_111000000000_000000100001_110100000001_000000000011_111000000000",	-- 4530
        b"100100110000_010000000000_010010100001_111000000000_000000000000_111000000000",	-- 4531
        b"010010000000_010011011000_000000100001_100011011110_100101100101_111011100000",	-- 4532
        b"110010000000_000100000000_000000100001_100011101110_100101100011_111000000000",	-- 4533
        b"100101101011_011000100001_010010100001_111110000000_000000000000_111000000000",	-- 4534
        b"010010001000_000000000000_000000100001_101110000000_000011100000_111000100000",	-- 4535
        b"110000100000_110000000000_000001111101_110011000010_100101100001_111000000000",	-- 4536
        b"010010001000_000000000000_000000100001_101110000000_000010010000_111000100000",	-- 4537
        b"010000110000_010011011000_000000100001_110011000001_100101100101_111000000000",	-- 4540
        b"010010001000_000000000000_000000100001_101110000000_000110000000_111000100000",	-- 4541
        b"010000110000_010011011000_000000100001_111110000000_000000000000_111000000000",	-- 4542
        b"010000110001_111011011000_001010100001_110001000001_100101111011_001001000000",	-- 4543
        b"110010000000_000000000000_000000100001_100011000001_100101100110_111000000000",	-- 4544
        b"010000110010_011011011000_001010100001_110001000001_100101111011_001001000000",	-- 4545
        b"110001101011_011000000000_000000100001_011110000000_000000000000_111000000000",	-- 4546
        b"110010000000_000000000000_000001011101_100001000011_001110010100_111000000000",	-- 4547
        b"010010001000_000000100000_000000100001_101110000000_111111111111_111000100000",	-- 4550
        b"100101101000_110000100000_011010100001_111110000000_000000000000_111000000000",	-- 4551
        b"010010001000_000000000000_000000100001_110011011111_100101101101_111000000000",	-- 4552
        b"010010001000_000000000000_000000100001_101110000000_000000000010_111000100000",	-- 4553
        b"010010000000_010000000000_000000100001_101110000000_000000000000_111011100000",	-- 4554
        b"010001101100_110000010000_000000100001_111110000000_000000000000_111000000000",	-- 4555
        b"100101101000_010000000000_010010100001_111110000000_000000000000_111000000000",	-- 4556
        b"100101101000_010000010000_010010100001_111110000000_000000000000_111000000000",	-- 4557
        b"100100110000_010000000000_010010100001_111110000000_000000000000_111000000000",	-- 4560
        b"010001101100_110000010000_000000100001_111110000000_000000000000_111000000000",	-- 4561
        b"010011000000_110000010000_000000100001_110100000001_000000000001_111000000000",	-- 4562
        b"100100110000_010000001000_000000100001_111000000000_000000000000_111000000000",	-- 4563
        b"110001101100_010000000001_111110100001_111110000000_000000000000_111000000000",	-- 4564
        b"100101101000_010000000000_010010100001_110100000001_000000000011_111000000000",	-- 4565
        b"100100110000_010000000000_010010100001_011000000000_000000000000_111000000000",	-- 4566
        b"110001101000_010000000000_000000110101_111010000011_000000000000_111010000000",	-- 4567
        b"110010000000_000000000000_000110100001_101110000000_000100100001_111000100000",	-- 4570
        b"010010000000_000100100000_000000100001_101010000001_000000000000_111010000000",	-- 4571
        b"010001101011_011011011000_001010100001_111110000000_000000000000_001001000000",	-- 4572
        b"110010000000_000000000000_000000100001_100001010001_100001101100_000000000000",	-- 4573
        b"010010000000_000100100000_000000100001_001110000000_000000000000_101001000000",	-- 4574
        b"110010000000_000000000000_000000100001_101010110001_000000000000_000000000000",	-- 4575
        b"110010000000_000000000000_000110100001_101110000000_000101011111_111000100000",	-- 4576
        b"110011000111_111000000000_000000100001_111110000000_000000000000_111010000000",	-- 4577
        b"110010000000_000000000000_000110100001_101110000000_000101100000_111000100000",	-- 4600
        b"110011000111_111000100000_000000100001_111110000000_000000000000_111010000000",	-- 4601
        b"010001101011_011000100000_000000100001_111110000000_000000000000_000000000000",	-- 4602
        b"100100110000_110000100000_010010100001_111110000000_000000000000_000000000000",	-- 4603
        b"010010000000_110000100000_000000100001_101110000000_000000000000_000011100000",	-- 4604
        b"011011000110_110000100000_000110100001_101110000000_000001010100_000000100000",	-- 4605
        b"010010000000_000000100000_000000100001_101110000000_000000000000_000010000000",	-- 4606
        b"011000111000_110000000000_001010100001_111110000000_000000000000_011001000000",	-- 4607
        b"010010000000_000000000000_000000100001_101110000000_000000000000_101001000000",	-- 4610
        b"010001101101_111000001000_000000100001_110011111001_100110001100_111000000000",	-- 4611
        b"010000110101_111000000000_000000100001_110011011011_100110001110_111000000000",	-- 4612
        b"010000110101_111000000000_000000100001_110011000001_100110100000_111000000000",	-- 4613
        b"010010001000_000000100000_000110100001_101110000000_000001101101_111000100000",	-- 4614
        b"110010000000_000000000000_000000100001_100011000001_100110100001_111000000000",	-- 4615
        b"010010001000_000000100000_000000100001_101110000000_110101101000_111000100000",	-- 4616
        b"100100110000_110000100000_010010100001_110001000001_100110101110_111000000000",	-- 4617
        b"011011000000_010000100000_000000100001_101110000000_000000000000_111000000000",	-- 4620
        b"010010001000_000000100000_000000100001_101110000000_100000001000_111000100000",	-- 4621
        b"100100110000_110000100000_010010100001_110001000001_100110101110_111000000000",	-- 4622
        b"110010111000_110000000000_000001101001_110011000011_100110100000_111000000000",	-- 4623
        b"110010000000_000000000000_000110100001_101110000000_000101101110_111000100000",	-- 4624
        b"011101101110_110000100010_000000100001_101110000000_000000000000_111010000000",	-- 4625
        b"011111111000_110000100000_000000100001_111110000000_000000000000_111010000000",	-- 4626
        b"010010000000_110000100000_000000100001_101110000000_000000000000_111011100000",	-- 4627
        b"110011001000_110000000000_000001101001_110011000010_100110011001_111000000000",	-- 4630
        b"010010001000_000000100000_000110100001_101110000000_000001110000_111000100000",	-- 4631
        b"110010000000_000000000000_000000100001_100001000001_100110101011_111000000000",	-- 4632
        b"110010000000_000000000000_000110100001_101110000000_000101011111_111000100000",	-- 4633
        b"010010000000_000000000000_000000100001_101110000000_000000000000_111010000000",	-- 4634
        b"110010000000_000000000000_000110100001_101110000000_000101100000_111000100000",	-- 4635
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 4636
        b"110001101100_110000000001_010110100001_111010000001_000000000000_111000000000",	-- 4637
        b"010010001000_000000100000_000110100001_101101000001_000001101010_111000100000",	-- 4640
        b"011001101000_110000000000_000110100001_101101000001_000001101000_111000100000",	-- 4641
        b"010010000000_000000100000_000000100001_101101000001_000000000000_111010000000",	-- 4642
        b"110001101000_110000000000_000001101001_110011000011_000000000000_111000100000",	-- 4643
        b"010011001111_111000100000_000110100001_110001000001_100110101001_111000000000",	-- 4644
        b"010010110101_111000000000_000000100001_101101000001_011111000000_111000100000",	-- 4645
        b"110011000111_110000000000_000001101001_111011000010_100111101010_111000000000",	-- 4646
        b"010010001000_000000000000_000000100001_101110000000_011110000000_111000100000",	-- 4647
        b"110010000000_000000000000_000000100001_101011000001_100111101010_111000000000",	-- 4650
        b"110010000000_000000000000_000000100001_001110000000_000000000000_111010000000",	-- 4651
        b"110010000000_000000000000_000001001001_101010000011_000000000000_111000000000",	-- 4652
        b"110011000111_111000000000_000000100001_110001000001_100110101111_111010000000",	-- 4653
        b"110011000111_111011011000_000000100001_110001000001_100110101111_111010000000",	-- 4654
        b"110011000111_111100100001_010110100001_111010000001_000000000000_111010000000",	-- 4655
        b"100100110000_110000100000_010010100001_111010000001_000000000000_111000000000",	-- 4656
        b"010001101000_110000100010_000110100001_111010000001_000000000000_111000000000",	-- 4657
        b"011101101100_010100010010_000000100001_110011011100_100110110010_111000000000",	-- 4660
        b"010011001111_111100000001_111110100001_110011000001_100110110011_111000000000",	-- 4661
        b"011111000110_111100000001_111110100001_110011000001_100110110011_111000000000",	-- 4662
        b"011111001111_010000000000_000000010100_000011111010_100110111111_111010000000",	-- 4663
        b"000110001000_000000100000_001010100001_101110000000_001111111110_111000100000",	-- 4664
        b"000101101000_110000100001_010010100001_111110000000_000000000000_111000000000",	-- 4665
        b"110011000000_010000100000_000001101001_110011000011_100111101101_111000000000",	-- 4666
        b"010011111000_010011011000_001010100001_110011011000_100110111011_001001000000",	-- 4667
        b"010011000110_111100000000_000000010100_110001000001_100100010110_111000000000",	-- 4670
        b"110010000000_000000000000_000000100001_100011000001_100110110010_111000000000",	-- 4671
        b"010001101100_010011011000_001010100001_111110000000_000000000000_001001000000",	-- 4672
        b"110010000000_000000000000_000000100001_100001010001_100001101100_000000000000",	-- 4673
        b"010010000000_000100100001_010110100001_001110000000_000000000000_101001000000",	-- 4674
        b"010001101100_110100100000_000000100001_111010110001_000000000000_000000000000",	-- 4675
        b"110010000000_000000000000_000000100001_100011000001_100101111110_000000000000",	-- 4676
        b"010001101100_010011011000_100110100001_110011010010_100110111010_111000000000",	-- 4677
        b"010010000000_000100100000_000000100001_101011010101_100111101001_111010000000",	-- 4700
        b"110010000000_000000000000_000000100001_100001010001_100001101100_111000000000",	-- 4701
        b"110001101100_110000000001_010110100001_111010000001_000000000000_111000000000",	-- 4702
        b"010001101011_011011011010_001010100001_110011000001_100111000101_010001000000",	-- 4703
        b"010001101011_011011011000_001010100001_111110000000_000000000000_010001000000",	-- 4704
        b"010001101100_110100100000_001010100001_011110000000_000000000000_101001000000",	-- 4705
        b"110010000000_000000000000_000000100001_101010110001_000000000000_000000000000",	-- 4706
        b"110010000000_000000000000_000000100001_100011000001_100101111110_000000000000",	-- 4707
        b"011101101100_010100000011_111110100001_110011000001_100111001010_111000000000",	-- 4710
        b"011111000110_111100000001_111110010110_110011100001_100111011111_111000000000",	-- 4711
        b"011011001111_010000000000_000000010110_000011111010_100111011111_111010000000",	-- 4712
        b"000110001000_000000100000_001010100001_101110000000_001111111110_111000100000",	-- 4713
        b"000101101000_110000100001_010010100001_111110000000_000000000000_111000000000",	-- 4714
        b"110011000000_010000100000_000001101001_110011000011_100111101101_111000000000",	-- 4715
        b"011011001110_111000000000_000110100001_101110000000_000100100011_111000100000",	-- 4716
        b"010010000000_000000100000_000000100001_101110000000_000000000000_111010000000",	-- 4717
        b"110010111000_110000000000_000001101001_110011000010_100111010100_111000000000",	-- 4720
        b"110010000000_000000000000_000110100001_101110000000_000001101001_111000100000",	-- 4721
        b"010010001000_000000100000_000000100001_101110000000_000000001000_111000100000",	-- 4722
        b"110011000111_111000100001_000000100001_111110000000_000000000000_111010000000",	-- 4723
        b"010011111000_010011011000_001010100001_110011011000_100111010111_010001000000",	-- 4724
        b"010011000110_111100000000_000000100001_110001000001_100100010100_111000000000",	-- 4725
        b"110010000000_000000000000_000000100001_100011000001_100111001001_111000000000",	-- 4726
        b"110010000000_000000000000_000000100001_100011101000_100111011100_000000000000",	-- 4727
        b"110011000100_111000000000_000000100001_010011100101_100111011010_111000000000",	-- 4730
        b"110010000000_000000000000_000001001001_100011000011_100111010101_111000000000",	-- 4731
        b"110010000000_000000000000_000000100001_100011000001_100111101110_111000000000",	-- 4732
        b"010001101100_010011011000_001010100001_111110000000_000000000000_010001000000",	-- 4733
        b"010001101100_110100100000_001010100001_011110000000_000000000000_101001000000",	-- 4734
        b"110010000000_000000000000_000000100001_101010110001_000000000000_000000000000",	-- 4735
        b"110010000000_000000000000_000000100001_100011000001_100101111110_000000000000",	-- 4736
        b"010001101100_010011011000_100110100001_110011010010_100111011011_111000000000",	-- 4737
        b"110010000000_000000000000_000000100001_101011010101_100111101001_111000000000",	-- 4740
        b"110011000111_111100100000_000000100001_111010000001_000000000000_111010000000",	-- 4741
        b"010010001000_000000000000_000000100001_101110000000_010001000000_111000100000",	-- 4742
        b"110010000000_000000000000_000000100001_101011000001_100111101010_111000000000",	-- 4743
        b"010010001000_000000000000_000000100001_111011000001_100111101110_111000000000",	-- 4744
        b"010010001000_000000000000_000000100001_101110000000_010000000000_111000100000",	-- 4745
        b"110010000000_000000000000_000000100001_101011000001_100111101010_111000000000",	-- 4746
        b"010010001000_000000000000_000000100001_101110000000_010100000000_111000100000",	-- 4747
        b"110010000000_000000000000_000000100001_101011000001_100111101010_111000000000",	-- 4750
        b"010010001000_000000000000_000000100001_101110000000_010111000000_111000100000",	-- 4751
        b"010010000000_010000000000_000000100001_100100000001_000000000010_111011100000",	-- 4752
        b"100100110000_010000000000_010010100001_111000000000_000000000000_111000000000",	-- 4753
        b"110010000000_000000000000_000000100001_100011000001_100111110011_111000000000",	-- 4754
        b"010000001000_000000000000_000000100001_110011000001_001001110110_111000000000",	-- 4755
        b"000110001000_000000100000_001010100001_101110000000_000000000001_111000100000",	-- 4756
        b"000101101000_110000100001_010010100001_111110000000_000000000000_111000000000",	-- 4757
        b"110011000000_010000100000_000001101001_110011000011_100111101101_111000000000",	-- 4760
        b"000101101100_111000100001_010010110101_110011000011_100111110011_111000000000",	-- 4761
        b"010011110000_110000000000_000000100001_111110000000_000000000000_111000000000",	-- 4762
        b"010010001000_000000100000_000000100001_101110000000_000000011111_111000100000",	-- 4763
        b"010010000000_110000100000_000000100001_101110000000_000000000000_111011100000",	-- 4764
        b"010011000000_110100001000_000000100001_110001100110_010100010100_111000000000",	-- 4765
        b"011010010110_111000000000_000110100001_101110000000_000001110100_111000100000",	-- 4766
        b"010011111100_010000000000_000000100001_111011100001_100111111010_111000000000",	-- 4767
        b"010010001000_000000100000_000000100001_101110000000_001000000000_111000100000",	-- 4770
        b"010010000000_110000100000_000000100001_100001000001_011001100000_111011100000",	-- 4771
        b"010001101000_010100100000_000000100001_110001011110_101000001010_111000000000",	-- 4772
        b"010010000000_000000100000_000000100001_001110000000_000000000000_111010000000",	-- 4773
        b"110001101000_110000000000_000001001001_110011000011_000000000000_111000100000",	-- 4774
        b"010010001000_000000000000_000000100001_101110000000_101000001100_111000100000",	-- 4775
        b"010000110111_111011110000_000000100001_110001000001_101000010001_111000000000",	-- 4776
        b"010010001000_000011011000_000000100001_101110000000_000101000000_111000100000",	-- 4777
        b"010000110010_011011011000_001010100001_110001000001_100111000100_010001000000",	-- 5000
        b"010001101000_011100100000_000000100001_110011100100_101000000011_111000000000",	-- 5001
        b"010001101011_110100110000_000000100001_110011000001_101000000101_111000000000",	-- 5002
        b"010001101011_011011011010_001010100001_110001000001_100111000100_010001000000",	-- 5003
        b"010001101011_110100100000_000000100001_111110000000_000000000000_111000000000",	-- 5004
        b"010001101011_011011011010_001010100001_110001000001_100111000100_010001000000",	-- 5005
        b"010001101011_011011011010_001010100001_110001000001_100101111011_001001000000",	-- 5006
        b"010010001000_000000000000_000000100001_110001000001_101000010001_111000000000",	-- 5007
        b"010001101100_110011100000_100000100001_110011100101_010011001101_111000000000",	-- 5010
        b"010010001000_000000011000_011000100001_110011000001_001100010000_111000000000",	-- 5011
        b"000110001000_000000000000_001010100001_101110000000_000000000000_111000100000",	-- 5012
        b"010011110000_010100100000_000000100001_111010000001_000000000000_111000000000",	-- 5013
        b"010010001000_000000000000_000000100001_101110000000_000000000100_111000100000",	-- 5014
        b"110010000000_000000000000_000000100001_101011000001_001001110110_111000000000",	-- 5015
        b"110010000000_000000000000_000000100001_100001000001_101000010001_111000000000",	-- 5016
        b"110010000000_000000000000_000110100001_101110000000_000001110100_111000100000",	-- 5017
        b"110011000111_111000000000_000000100001_111010000001_000000000000_111010000000",	-- 5020
        b"110010000000_000000000000_000110100001_101110000000_000001101000_111000100000",	-- 5021
        b"110001101000_010000000000_000000100001_111010000001_000000000000_111010000000",	-- 5022
    );
micro2: Note: Dump of DROM Statements.
width = 96
    constant DROM : DROM_t := (
        --000000000011_111111112222_222222333333_333344444444_445555555555_666666666677_777777778888_888888999999
        --012345678901_234567890123_456789012345_678901234567_890123456789_012345678901_234567890123_456789012345
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011000111110_001011000100",	-- 0000
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0001
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0002
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0003
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011001000000_001011000100",	-- 0004
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011001100001_001011000100",	-- 0005
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011001101001_001011000100",	-- 0006
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011001101011_001011000100",	-- 0007
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0010
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0011
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0012
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0013
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011001101101_001011000100",	-- 0014
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011010101111_001011000100",	-- 0015
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011010111101_001011000100",	-- 0016
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011011000000_001011000100",	-- 0017
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0020
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011011101110_001011000100",	-- 0021
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011100001010_001011000100",	-- 0022
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011011011011_001011000100",	-- 0023
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011011000011_001011000100",	-- 0024
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_011011010110_001011000100",	-- 0025
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0026
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0027
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0030
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0031
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0032
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0033
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0034
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0035
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0036
        b"010101001000_001011000100_001110000000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0037
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011011111010_001011000100",	-- 0040
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100001000_001011000100",	-- 0041
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100000011_001011000100",	-- 0042
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011011111110_001011000100",	-- 0043
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100001111_001011000100",	-- 0044
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100100001_001011000100",	-- 0045
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100101101_001011000100",	-- 0046
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0047
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011011111000_001011000100",	-- 0050
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100000101_001011000100",	-- 0051
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100000000_001011000100",	-- 0052
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011011111011_001011000100",	-- 0053
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100011100_001011000100",	-- 0054
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100100100_001011000100",	-- 0055
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_011100101010_001011000100",	-- 0056
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0057
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0060
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0061
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0062
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0063
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0064
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0065
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0066
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0067
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0070
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0071
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0072
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0073
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0074
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0075
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0076
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0077
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0100
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0101
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0102
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0103
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0104
        b"001101010110_010101001000_010100101101_010100110001_001011000100_001011000100_001110011111_001011000100",	-- 0105
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0106
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0107
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0110
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0111
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0112
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0113
        b"001100111100_010001110011_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0114
        b"001100111100_010001111010_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0115
        b"001100111100_010001111101_100100001010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0116
        b"001100111100_010001111101_100100001010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0117
        b"001100111110_100011100101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0120
        b"001100111110_001110110110_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0121
        b"001101001001_010000100000_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0122
        b"010111101000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0123
        b"001100111010_100011111111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0124
        b"001100111010_001110110110_100011111111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0125
        b"001101001001_010000100000_010000101101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0126
        b"001101001001_010000110001_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0127
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0130
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0131
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0132
        b"001101001000_001111011001_100001010111_001110111101_001011000100_001011000100_001110011111_001011000100",	-- 0133
        b"001101001110_001111110000_010000001000_010000001001_001011000100_001011000100_001110011111_001011000100",	-- 0134
        b"001101001001_001111011010_001011000100_010000001001_001011000100_001011000100_001110011111_001011000100",	-- 0135
        b"001101001101_001111110000_010000001000_010000010001_001011000100_001011000100_001110011111_001011000100",	-- 0136
        b"001101001000_001111011010_001011000100_010000010001_001011000100_001011000100_001110011111_001011000100",	-- 0137
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0140
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0141
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0142
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0143
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0144
        b"001101010110_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0145
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0146
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0147
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0150
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0151
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0152
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0153
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0154
        b"001101010110_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0155
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0156
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0157
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0160
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0161
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0162
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0163
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0164
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0165
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0166
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0167
        b"001101001001_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0170
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0171
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0172
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0173
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0174
        b"001101001000_010000110001_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0175
        b"001101001101_010000110001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0176
        b"001101001101_010000110001_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0177
        b"001101001001_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0200
        b"010000110001_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0201
        b"001101011001_100011111001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0202
        b"001101001110_100011101010_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0203
        b"001101001001_010000110100_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0204
        b"010000110010_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0205
        b"001101011001_010000110100_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0206
        b"001101001101_010000110100_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0207
        b"001101001001_010000110110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0210
        b"001101010111_010000110110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0211
        b"001101011010_010000110110_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0212
        b"001101001110_010000110110_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0213
        b"001101001001_010000110101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0214
        b"010000110001_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0215
        b"001101011010_010000110101_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0216
        b"001101001110_010000110101_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0217
        b"001101001000_010001000011_010001001100_100011100010_001011000100_001011000100_001110011111_001011000100",	-- 0220
        b"001101010110_010001000011_010001001100_100011100010_001011000100_001011000100_001110011111_001011000100",	-- 0221
        b"001101001101_010001000011_010001001100_100011110011_001011000100_001011000100_001110011111_001011000100",	-- 0222
        b"001101001101_010001000011_010001001100_100011101111_001011000100_001011000100_001110011111_001011000100",	-- 0223
        b"001101001000_010001000011_100011100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0224
        b"001101010110_010001000011_100011100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0225
        b"001101001101_010001000011_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0226
        b"001101001101_010001000011_100011011100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0227
        b"001101001000_010001001111_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0230
        b"001101010110_010001001111_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0231
        b"001101001101_010001001111_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0232
        b"001101001101_010001001111_100011011100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0233
        b"001101001000_010001010010_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0234
        b"001101010110_010001010010_100011100000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0235
        b"001101001101_010001010010_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0236
        b"001101001101_010001010010_100011011100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0237
        b"001101011010_010010000001_010010001000_010010001100_001011000100_001011000100_001110011111_001011000100",	-- 0240
        b"001101011001_010010000001_010010100001_010010100011_001011000100_001011000100_001110011111_001011000100",	-- 0241
        b"001101011001_010010000001_010010011001_010010011011_001011000100_001011000100_001110011111_001011000100",	-- 0242
        b"001101011010_010011111010_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0243
        b"001100111010_010001111110_010010001110_010010010110_001011000100_001011000100_001110011111_001011000100",	-- 0244
        b"001100111010_010010000000_010010100101_010010100111_001011000100_001011000100_001110011111_001011000100",	-- 0245
        b"001100111010_010010000000_010010011101_010010011111_001011000100_001011000100_001110011111_001011000100",	-- 0246
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0247
        b"001101001101_100011110001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0250
        b"001101011001_010010101001_010010111100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0251
        b"001101011001_010011000000_010110101000_100011100010_001011000100_001011000100_001110011111_001011000100",	-- 0252
        b"001101011001_010011000000_010110100001_100011100010_001011000100_001011000100_001110011111_001011000100",	-- 0253
        b"010011000010_001011000100_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0254
        b"010100000000_001011000100_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0255
        b"001101001001_010100000110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0256
        b"010100100101_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0257
        b"001101011001_010101001000_010100110110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0260
        b"001101001000_010101001001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0261
        b"001101011001_010101001000_010101011000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0262
        b"001101011001_010101001000_010101110001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0263
        b"010101001000_010101111111_010101111011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0264
        b"010101001000_010110000100_010101111011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0265
        b"001101011001_010110000101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0266
        b"001101011001_010110001010_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0267
        b"001101001000_010000111011_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0270
        b"001101010110_010000111011_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0271
        b"001101001101_010000111011_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0272
        b"001101001101_010000111011_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0273
        b"001101001000_010000111110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0274
        b"001101010110_010000111110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0275
        b"001101001101_010000111110_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0276
        b"001101001101_010000111110_100011101111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0277
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0300
        b"001101010110_010110001110_010110010101_001100010000_001011000100_001011000100_001110011111_010110100111",	-- 0301
        b"001101010110_010110001110_010110010111_001100010000_001011000100_001011000100_001110011111_010011000101",	-- 0302
        b"001101010110_010110001110_010110011001_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0303
        b"001101010110_010110001110_010110011010_001100010000_001011000100_001011000100_001110011111_010011010011",	-- 0304
        b"001101010110_010110001110_010110011011_001100010000_001011000100_001011000100_001110011111_010011010110",	-- 0305
        b"001101010110_010110001110_010110011101_001100010000_001011000100_001011000100_001110011111_010011011100",	-- 0306
        b"001101010110_010110001110_010110011111_001100010000_001011000100_001011000100_001110011111_010011100001",	-- 0307
        b"001101001001_001100010000_001011000100_001011000100_001011000100_001011000100_001110011111_010011101000",	-- 0310
        b"001101001000_010110001110_010110010101_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0311
        b"001101001000_010110001110_010110010111_001100010000_001011000100_001011000100_001110011111_010011101010",	-- 0312
        b"001101001000_010110001110_010110011001_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0313
        b"001101001000_010110001110_010110011010_001100010000_001011000100_001011000100_001110011111_010011110111",	-- 0314
        b"001101001000_010110001110_010110011011_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0315
        b"001101001000_010110001110_010110011101_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0316
        b"001101001000_010110001110_010110011111_001100010000_001011000100_001011000100_001110011111_001110011111",	-- 0317
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0320
        b"001101011010_010110100001_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0321
        b"001101011010_010110100011_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0322
        b"001101011010_010110100101_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0323
        b"010110100111_001011000100_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0324
        b"001101011010_010110101000_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0325
        b"001101011010_010110101010_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0326
        b"001101011010_010110101100_001011000100_001100010000_001011000100_001011000100_001110011111_001011000100",	-- 0327
        b"001101001001_010110101110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0330
        b"001101001001_010110010101_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0331
        b"001101001001_010110010111_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0332
        b"001101001001_010110011001_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0333
        b"001101001001_010110011010_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0334
        b"001101001001_010110011011_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0335
        b"001101001001_010110011101_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0336
        b"001101001001_010110011111_001011000100_010110101110_001011000100_001011000100_001110011111_001011000100",	-- 0337
        b"001101011001_010110001111_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0340
        b"001101011001_010110001111_010110100001_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0341
        b"001101011001_010110001111_010110100011_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0342
        b"001101011001_010110001111_010110100101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0343
        b"001101011001_010110001111_010110100111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0344
        b"001101011001_010110001111_010110101000_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0345
        b"001101011001_010110001111_010110101010_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0346
        b"001101011001_010110001111_010110101100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0347
        b"001101001110_010110001111_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0350
        b"001101001110_010110001111_010110010101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0351
        b"001101001110_010110001111_010110010111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0352
        b"001101001110_010110001111_010110011001_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0353
        b"001101001110_010110001111_010110011010_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0354
        b"001101001110_010110001111_010110011011_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0355
        b"001101001110_010110001111_010110011101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0356
        b"001101001110_010110001111_010110011111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0357
        b"001101011001_010110010010_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0360
        b"001101011001_010110010010_010110100001_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0361
        b"001101011001_010110010010_010110100011_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0362
        b"001101011001_010110010010_010110100101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0363
        b"001101011001_010110010010_010110100111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0364
        b"001101011001_010110010010_010110101000_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0365
        b"001101011001_010110010010_010110101010_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0366
        b"001101011001_010110010010_010110101100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0367
        b"001101001110_010110010010_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0370
        b"001101001110_010110010010_010110010101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0371
        b"001101001110_010110010010_010110010111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0372
        b"001101001110_010110010010_010110011001_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0373
        b"001101001110_010110010010_010110011010_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0374
        b"001101001110_010110010010_010110011011_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0375
        b"001101001110_010110010010_010110011101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0376
        b"001101001110_010110010010_010110011111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0377
        b"010110110000_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0400
        b"010110110000_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0401
        b"010110110000_100011111001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0402
        b"010110110000_100011110000_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0403
        b"001101001000_010110110001_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0404
        b"001101010110_010110110001_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0405
        b"001101001101_010110110001_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0406
        b"001101001101_010110110001_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0407
        b"001101001000_010110110010_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0410
        b"001101010110_010110110010_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0411
        b"001101001101_010110110010_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0412
        b"001101001101_010110110010_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0413
        b"001101001001_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0414
        b"010110110011_001011000100_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0415
        b"001101001110_100011110011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0416
        b"001101001110_100011110000_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0417
        b"001101001000_010110110101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0420
        b"001101010110_010110110101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0421
        b"001101001101_010110110101_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0422
        b"001101001101_010110110101_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0423
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0424
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0425
        b"001101011001_100011111001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0426
        b"001101011001_100011111001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0427
        b"001101001000_010110110110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0430
        b"001101010110_010110110110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0431
        b"001101001101_010110110110_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0432
        b"001101001101_010110110110_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0433
        b"001101001000_010110111000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0434
        b"001101010110_010110111000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0435
        b"001101001101_010110111000_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0436
        b"001101001101_010110111000_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0437
        b"001101001000_010110111001_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0440
        b"001101010110_010110111001_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0441
        b"001101001101_010110111001_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0442
        b"001101001101_010110111001_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0443
        b"001101001000_010110111011_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0444
        b"001101010110_010110111011_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0445
        b"001101001101_010110111011_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0446
        b"001101001101_010110111011_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0447
        b"001101011001_010110111100_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0450
        b"001101011001_010110111100_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0451
        b"001101011001_010110111100_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0452
        b"001101011001_010110111100_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0453
        b"001101001000_010110111101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0454
        b"001101010110_010110111101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0455
        b"001101001101_010110111101_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0456
        b"001101001101_010110111101_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0457
        b"001101001001_010110111110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0460
        b"001101010111_010110111110_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0461
        b"001101001110_010110111110_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0462
        b"001101001110_010110111110_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0463
        b"001101001000_010110111111_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0464
        b"001101010110_010110111111_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0465
        b"001101001101_010110111111_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0466
        b"001101001101_010110111111_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0467
        b"001101001000_010111000000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0470
        b"001101010110_010111000000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0471
        b"001101001101_010111000000_100011110011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0472
        b"001101001101_010111000000_100011110000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0473
        b"010111000001_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0474
        b"010111000001_100011100011_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0475
        b"010111000001_100011111001_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0476
        b"010111000001_100011110000_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0477
        b"001101001000_010111000010_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0500
        b"001101011001_010111000011_100011100010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0501
        b"001101001101_010111001001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0502
        b"001101001110_100011101010_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0503
        b"001101001000_010111001010_100011101000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0504
        b"001101010110_010111001010_100011101000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0505
        b"001101001101_010111001000_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0506
        b"001101001101_010111001011_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0507
        b"001101001001_010111001100_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0510
        b"001101010111_010111001100_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0511
        b"001101011001_010111001100_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0512
        b"001101001110_010111001100_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0513
        b"001101001001_010000110100_010111001100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0514
        b"010000110010_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0515
        b"001101011001_010000110100_010111001100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0516
        b"001101001110_010000110100_010111001100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0517
        b"001101001001_010111001111_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0520
        b"001101010111_010111001111_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0521
        b"001101011001_010111001111_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0522
        b"001101001110_010111001111_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0523
        b"001101001001_010000110100_010111001111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0524
        b"001101010111_010000110100_010111001111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0525
        b"001101011001_010000110100_010111001111_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0526
        b"001101001110_010000110100_010111001111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0527
        b"001101001001_010111001110_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0530
        b"001101010111_010111001110_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0531
        b"001101011010_010111001110_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0532
        b"001101001110_010111001110_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0533
        b"001101001001_010000110100_010111001101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0534
        b"001101010111_010000110100_010111001101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0535
        b"001101011010_010000110100_010111001101_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0536
        b"001101001110_010000110100_010111001101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0537
        b"001101001000_010111010000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0540
        b"001101010110_010111010000_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0541
        b"001101001101_010111010010_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0542
        b"001101001110_100011101010_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0543
        b"001101001000_010111010011_100011101000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0544
        b"001101010110_010111010011_100011101000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0545
        b"001101001101_010111010001_100011111001_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0546
        b"001101001101_010111010100_100011101010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0547
        b"001101001001_010111010101_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0550
        b"010000110001_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0551
        b"001101011001_010111010101_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0552
        b"001101001110_010111010101_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0553
        b"001101001001_010000110100_010111010101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0554
        b"001101010111_010000110100_010111010101_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0555
        b"001101011001_010000110100_010111010101_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0556
        b"001101001110_010000110100_010111010101_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0557
        b"001101001001_010111010111_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0560
        b"001101010111_010111010111_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0561
        b"001101011001_010111010111_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0562
        b"001101001110_010111010111_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0563
        b"001101001001_010000110100_010111010111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0564
        b"001101010111_010000110100_010111010111_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0565
        b"001101011001_010000110100_010111010111_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0566
        b"001101001110_010000110100_010111010111_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0567
        b"001101001001_010111010110_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0570
        b"001101010111_010111010110_001011000100_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0571
        b"001101011010_010111010110_001011000100_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0572
        b"001101001110_010111010110_001011000100_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0573
        b"001101001001_010000110100_010111010110_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0574
        b"001101010111_010000110100_010111010110_100011100011_001011000100_001011000100_001110011111_001011000100",	-- 0575
        b"001101011010_010000110100_010111010110_100011111001_001011000100_001011000100_001110011111_001011000100",	-- 0576
        b"001101001110_010000110100_010111010110_100011101010_001011000100_001011000100_001110011111_001011000100",	-- 0577
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0600
        b"100001010111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0601
        b"010111011000_010111100001_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0602
        b"010111011001_010111100001_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0603
        b"010111011000_010111100010_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0604
        b"010111011001_010111100010_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0605
        b"010111011000_010111100011_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0606
        b"010111011001_010111100011_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0607
        b"010111011011_001100010000_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0610
        b"010111011110_001100010000_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0611
        b"010111011011_010111100001_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0612
        b"010111011110_010111100001_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0613
        b"010111011011_010111100010_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0614
        b"010111011110_010111100010_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0615
        b"010111011011_010111100011_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0616
        b"010111011110_010111100011_001100010000_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0617
        b"010111011000_010111100101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0620
        b"010111011001_010111100101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0621
        b"010111011000_010111100001_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0622
        b"010111011001_010111100001_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0623
        b"010111011000_010111100010_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0624
        b"010111011001_010111100010_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0625
        b"010111011000_010111100011_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0626
        b"010111011001_010111100011_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0627
        b"010111011011_010111100101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0630
        b"010111011110_010111100101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0631
        b"010111011011_010111100001_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0632
        b"010111011110_010111100001_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0633
        b"010111011011_010111100010_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0634
        b"010111011110_010111100010_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0635
        b"010111011011_010111100011_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0636
        b"010111011110_010111100011_010111100101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0637
        b"010111011000_010111100110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0640
        b"010111011001_010111100110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0641
        b"010111011000_010111100001_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0642
        b"010111011001_010111100001_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0643
        b"010111011000_010111100010_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0644
        b"010111011001_010111100010_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0645
        b"010111011000_010111100011_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0646
        b"010111011001_010111100011_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0647
        b"010111011011_010111100110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0650
        b"010111011110_010111100110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0651
        b"010111011011_010111100001_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0652
        b"010111011110_010111100001_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0653
        b"010111011011_010111100010_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0654
        b"010111011110_010111100010_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0655
        b"010111011011_010111100011_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0656
        b"010111011110_010111100011_010111100110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0657
        b"010111011000_010111100111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0660
        b"010111011001_010111100111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0661
        b"010111011000_010111100001_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0662
        b"010111011001_010111100001_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0663
        b"010111011000_010111100010_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0664
        b"010111011001_010111100010_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0665
        b"010111011000_010111100011_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0666
        b"010111011001_010111100011_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0667
        b"010111011011_010111100111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0670
        b"010111011110_010111100111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0671
        b"010111011011_010111100001_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0672
        b"010111011110_010111100001_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0673
        b"010111011011_010111100010_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0674
        b"010111011110_010111100010_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0675
        b"010111011011_010111100011_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0676
        b"010111011110_010111100011_010111100111_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0677
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0700
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0701
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0702
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0703
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0704
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0705
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0706
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0707
        b"100000011000_001101011100_100000011010_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0710
        b"100000011000_001101011100_100000011100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0711
        b"100000011000_001101011101_100011100011_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0712
        b"100000011000_100000011110_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0713
        b"100000011000_001101011100_100001010101_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0714
        b"100000011000_001101011100_100001010110_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0715
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0716
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0717
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0720
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0721
        b"011100101111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0722
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0723
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0724
        b"001110011111_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0725
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0726
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0727
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0730
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0731
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0732
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0733
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0734
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0735
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0736
        b"011000110100_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0737
        b"010111101010_010111111101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0740
        b"010111101010_011000000101_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0741
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0742
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0743
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0744
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0745
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0746
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0747
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0750
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0751
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0752
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0753
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0754
        b"010111101010_011000001111_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0755
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0756
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0757
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0760
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0761
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0762
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0763
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0764
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0765
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0766
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0767
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0770
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0771
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0772
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0773
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0774
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0775
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0776
        b"011000111000_001011000100_001011000100_001011000100_001011000100_001011000100_001110011111_001011000100",	-- 0777
    );
